magic
tech sky130A
magscale 1 2
timestamp 1743030000
<< checkpaint >>
rect 0 0 8944 6440
use JNWTR_RPPO2 x5 ../JNW_TR_SKY130A
transform 1 0 0 0 1 0
box 0 0 1448 3440
use JNWTR_RPPO16 x6 ../JNW_TR_SKY130A
transform 1 0 2128 0 1 0
box 2128 0 6600 3440
use JNWATR_PCH_12C5F0 xb1 ../JNW_ATR_SKY130A
transform 1 0 7280 0 1 0
box 7280 0 8944 800
use JNWATR_PCH_12C5F0 xb2 ../JNW_ATR_SKY130A
transform 1 0 7280 0 1 800
box 7280 800 8944 1600
use JNWATR_PCH_4C1F2 xli1 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 4040
box 0 4040 1152 4840
use JNWATR_NCH_4C5F0 xlo1 ../JNW_ATR_SKY130A
transform 1 0 1832 0 1 4040
box 1832 4040 2984 4840
use JNWATR_PCH_4C5F0 xlo2 ../JNW_ATR_SKY130A
transform 1 0 1832 0 1 4840
box 1832 4840 2984 5640
use JNWATR_NCH_4C5F0 xlo3 ../JNW_ATR_SKY130A
transform 1 0 1832 0 1 5640
box 1832 5640 2984 6440
use JNWATR_NCH_4C5F0 xri1 ../JNW_ATR_SKY130A
transform 1 0 3664 0 1 4040
box 3664 4040 4816 4840
use JNWATR_PCH_4C1F2 xri2 ../JNW_ATR_SKY130A
transform 1 0 3664 0 1 4840
box 3664 4840 4816 5640
use JNWATR_NCH_4C5F0 xro1 ../JNW_ATR_SKY130A
transform 1 0 5496 0 1 4040
box 5496 4040 6648 4840
use JNWATR_PCH_4C5F0 xro2 ../JNW_ATR_SKY130A
transform 1 0 5496 0 1 4840
box 5496 4840 6648 5640
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 8944 6440
<< end >>
