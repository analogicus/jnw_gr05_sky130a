magic
tech sky130A
magscale 1 2
timestamp 1744566877
<< locali >>
rect -10229 7451 -2855 7452
rect -10229 7187 1768 7451
rect -10229 5057 -9964 7187
rect -11437 4902 -9964 5057
rect -5585 4954 1768 7187
rect -11437 4066 -11282 4902
rect -10387 4066 -10232 4902
rect -11437 4061 -10232 4066
rect -10229 4104 -9964 4902
rect -5628 4928 1768 4954
rect -9563 4180 -9396 4420
rect -6172 4180 -5991 4420
rect -5628 4104 -3697 4928
rect -10229 4061 -3697 4104
rect -11437 4027 -3697 4061
rect -3081 4310 1768 4928
rect -3081 4027 -1583 4310
rect -11437 3989 -1583 4027
rect -11437 3928 -10232 3989
rect -10229 3928 -1583 3989
rect -11473 3887 -1583 3928
rect -11475 3839 -1583 3887
rect -11475 3637 -8051 3839
rect -11469 3459 -8051 3637
rect -7872 3480 -1583 3839
rect -525 4212 1768 4310
rect -525 3480 926 4212
rect -7872 3459 926 3480
rect -11469 2646 -11280 3459
rect -10416 3330 -10061 3459
rect -10416 3008 -10040 3330
rect -10421 2646 -10040 3008
rect -9985 2686 -9846 3459
rect -8990 3388 -8487 3459
rect -8990 2690 -8851 3388
rect -9985 2646 -9839 2686
rect -9021 2646 -8851 2690
rect -8815 2661 -8487 3388
rect -7614 3207 926 3459
rect 1576 3207 1768 3380
rect -7614 3140 1768 3207
rect -7614 2673 -7425 3140
rect -8815 2646 -8439 2661
rect -7621 2646 -7425 2673
rect -7420 2646 -7279 3140
rect -6896 2942 -6444 2948
rect -6896 2762 -6890 2942
rect -6710 2762 -6444 2942
rect -6896 2756 -6444 2762
rect -11469 2627 -7279 2646
rect -11405 2458 -7279 2627
rect -11473 2108 -7279 2458
rect -11473 2079 -7754 2108
rect -11474 1303 -11262 2031
rect -10421 1876 -9839 2031
rect -11474 1257 -11239 1303
rect -10421 1261 -9876 1876
rect -9021 1445 -8439 2079
rect -7621 1782 -7425 2108
rect -9021 1261 -8474 1445
rect -10421 1260 -8243 1261
rect -7614 1260 -7425 1782
rect -10421 1257 -7425 1260
rect -11474 1183 -7425 1257
rect -11474 1125 -7465 1183
rect -7420 1125 -7279 2108
rect -11474 1071 -7279 1125
rect -11474 1068 -9937 1071
rect -11474 1058 -11239 1068
rect -11474 1027 -11162 1058
rect -10285 1027 -9937 1068
rect -9015 1027 -7279 1071
rect -11474 858 -7279 1027
rect -11476 823 -7279 858
rect -11476 792 -7268 823
rect -11476 746 -10942 792
rect -11474 -461 -10982 746
rect -7773 -51 -7268 792
rect -5895 79 -4640 3140
rect -1465 3015 1768 3140
rect -1465 3012 925 3015
rect -1465 2180 -915 3012
rect -2172 1940 773 2180
rect -2172 1840 538 1940
rect -3612 737 -3420 880
rect -2463 737 -2172 752
rect -3612 688 -2172 737
rect -1466 688 538 1840
rect -3612 380 538 688
rect -2463 318 538 380
rect -5876 -51 -4640 79
rect -7773 -140 -4640 -51
rect -7773 -444 -5046 -140
rect -5010 -268 -4640 -140
rect -4281 -268 -4089 -6
rect -7790 -461 -5036 -444
rect -11474 -556 -5036 -461
rect -11474 -770 -5094 -556
rect -11474 -4974 -10982 -770
rect -7773 -902 -5094 -770
rect -11480 -5106 -10982 -4974
rect -7717 -2084 -5094 -902
rect -1466 -852 538 318
rect -1466 -1032 -628 -852
rect -436 -1032 538 -852
rect -1466 -1358 538 -1032
rect -2058 -1550 538 -1358
rect -7717 -2276 -4990 -2084
rect -7717 -5106 -7408 -2276
rect -1759 -2513 538 -1550
rect -1670 -2527 538 -2513
rect -1670 -2693 539 -2527
rect -1862 -2719 539 -2693
rect -1862 -2978 -1670 -2719
rect -1754 -2996 -1734 -2978
rect -1810 -3188 -1734 -2996
rect -664 -3188 -604 -3060
rect -172 -3188 543 -3060
rect -1862 -3642 -1734 -3494
rect 351 -3636 543 -3188
rect -129 -3642 543 -3636
rect -1862 -3686 -845 -3642
rect -1111 -3822 -845 -3686
rect -129 -3822 -123 -3642
rect 57 -3670 543 -3642
rect 57 -3822 223 -3670
rect -1111 -4020 -667 -3822
rect -129 -3828 223 -3822
rect 100 -3850 223 -3828
rect 415 -3850 543 -3670
rect 100 -4020 543 -3850
rect -1111 -4212 543 -4020
rect -11480 -5178 -7408 -5106
rect -11480 -5370 -6534 -5178
<< viali >>
rect -9791 4180 -9563 4420
rect -5991 4180 -5763 4420
rect -6890 2762 -6710 2942
rect -6444 2756 -6264 2948
rect -4281 -6 -4089 174
rect -628 -1032 -436 -852
rect -1862 -2693 -1670 -2513
rect -845 -3822 -665 -3642
rect -123 -3822 57 -3642
rect 223 -3850 415 -3670
<< metal1 >>
rect -9797 4420 -9557 4432
rect -10984 4180 -9791 4420
rect -9563 4180 -9557 4420
rect -6001 4420 -2564 4504
rect -6001 4312 -5991 4420
rect -9797 4168 -9557 4180
rect -5997 4180 -5991 4312
rect -5763 4312 -2564 4420
rect -5763 4180 -4516 4312
rect -5997 4168 -5757 4180
rect -3397 3672 -2434 3864
rect -2311 3862 -960 3864
rect -2311 3672 -1929 3862
rect -1935 3670 -1929 3672
rect -1737 3672 -960 3862
rect -1737 3670 -1731 3672
rect -3387 3606 -1535 3608
rect -3387 3544 -1164 3606
rect -1599 3542 -1164 3544
rect -1599 3444 -1535 3542
rect -1604 3381 -1535 3444
rect -10859 2900 -9478 3092
rect -6450 2948 -6258 2960
rect -10859 1648 -10667 2900
rect -9670 1648 -9478 2900
rect -7896 2942 -6444 2948
rect -7896 2762 -6890 2942
rect -6710 2762 -6444 2942
rect -7896 2756 -6444 2762
rect -6264 2756 -3304 2948
rect -3096 2756 -2404 2948
rect -6450 2744 -6258 2756
rect -4558 1863 -4494 2756
rect -1604 2564 -1540 3381
rect 1480 2820 1672 2844
rect -418 2628 264 2820
rect 398 2628 1672 2820
rect -2276 2372 -1929 2564
rect -1737 2372 -492 2564
rect -446 2372 388 2564
rect -1604 2308 -1540 2372
rect 1480 2308 1672 2628
rect -2932 2244 -768 2308
rect -202 2244 126 2308
rect 553 2244 1672 2308
rect -4564 1799 -4558 1863
rect -4494 1799 -4488 1863
rect -10859 1456 -3260 1648
rect -2999 1456 -2540 1648
rect -4558 1245 -4494 1251
rect -4558 58 -4494 1181
rect -4281 832 -4089 838
rect -4281 180 -4089 640
rect -4293 174 -4077 180
rect -4293 -6 -4281 174
rect -4089 -6 -4077 174
rect -3900 114 -3836 1456
rect -2304 1261 -1740 1264
rect -2304 1072 -1929 1261
rect -1935 1069 -1929 1072
rect -1737 1069 -1731 1261
rect -1604 1008 -1540 2244
rect -3042 944 -1532 1008
rect -3414 557 -3284 749
rect -3900 62 -2758 114
rect -3900 50 -2694 62
rect -4293 -12 -4077 -6
rect -640 -852 -424 -846
rect -640 -1032 -628 -852
rect -436 -1032 -424 -852
rect -640 -1038 -424 -1032
rect -628 -1133 -436 -1038
rect -628 -1331 -436 -1325
rect -1862 -2210 -1670 -2204
rect -1862 -2507 -1670 -2402
rect -1874 -2513 -1658 -2507
rect -1874 -2693 -1862 -2513
rect -1670 -2693 -1658 -2513
rect -1874 -2699 -1658 -2693
rect -664 -3380 -478 -3374
rect 1480 -3380 1672 2244
rect -664 -3572 -478 -3566
rect -318 -3572 1672 -3380
rect -857 -3642 69 -3636
rect -857 -3822 -845 -3642
rect -665 -3822 -123 -3642
rect 57 -3822 69 -3642
rect -857 -3828 69 -3822
rect 211 -3670 427 -3664
rect 211 -3850 223 -3670
rect 415 -3850 427 -3670
rect 211 -3856 427 -3850
rect -1282 -3956 -550 -3892
rect 223 -3909 415 -3856
rect 223 -4107 415 -4101
<< via1 >>
rect -1929 3670 -1737 3862
rect -1929 2372 -1737 2564
rect -4558 1799 -4494 1863
rect -4558 1181 -4494 1245
rect -4281 640 -4089 832
rect -1929 1069 -1737 1261
rect -628 -1325 -436 -1133
rect -1862 -2402 -1670 -2210
rect -664 -3566 -478 -3380
rect 223 -4101 415 -3909
<< metal2 >>
rect -1929 3862 -1737 3868
rect -1929 2564 -1737 3670
rect -4558 1863 -4494 1869
rect -4558 1245 -4494 1799
rect -1929 1261 -1737 2372
rect -4564 1181 -4558 1245
rect -4494 1181 -4488 1245
rect -1929 832 -1737 1069
rect -4287 640 -4281 832
rect -4089 640 -1737 832
rect -634 -1325 -628 -1133
rect -436 -1325 -430 -1133
rect -628 -1388 -436 -1325
rect -628 -1579 -436 -1570
rect -1868 -2402 -1862 -2210
rect -1670 -2402 -1583 -2210
rect -1401 -2402 -1392 -2210
rect -1014 -3572 -1005 -3380
rect -823 -3566 -664 -3380
rect -478 -3566 -262 -3380
rect -86 -3566 -77 -3380
rect -823 -3572 -637 -3566
rect 217 -4101 223 -3909
rect 415 -4101 421 -3909
rect 223 -4151 415 -4101
rect 223 -4342 415 -4333
<< via2 >>
rect -628 -1570 -436 -1388
rect -1583 -2402 -1401 -2210
rect -1005 -3572 -823 -3380
rect -262 -3566 -86 -3380
rect 223 -4333 415 -4151
<< metal3 >>
rect -633 -1388 -431 -1383
rect -633 -1570 -628 -1388
rect -436 -1570 -431 -1388
rect -633 -1575 -431 -1570
rect -628 -1624 -436 -1575
rect -628 -1820 -436 -1814
rect -1588 -2210 -1396 -2205
rect -1588 -2402 -1583 -2210
rect -1401 -2402 -1387 -2210
rect -1197 -2402 -1191 -2210
rect -1588 -2407 -1396 -2402
rect -1010 -3380 -818 -2752
rect -1010 -3572 -1005 -3380
rect -823 -3572 -818 -3380
rect -1010 -4017 -818 -3572
rect -267 -3380 -81 -2782
rect -267 -3566 -262 -3380
rect -86 -3566 -81 -3380
rect -267 -4089 -81 -3566
rect 218 -4151 420 -4146
rect 218 -4333 223 -4151
rect 415 -4333 420 -4151
rect 218 -4338 420 -4333
rect 223 -4446 415 -4338
rect 223 -4642 415 -4636
<< via3 >>
rect -628 -1814 -436 -1624
rect -1387 -2402 -1197 -2210
rect 223 -4636 415 -4446
<< metal4 >>
rect -629 -1624 -435 -1623
rect -629 -1814 -628 -1624
rect -436 -1814 -435 -1624
rect -629 -1815 -435 -1814
rect -1388 -2210 -1196 -2209
rect -1388 -2402 -1387 -2210
rect -1197 -2402 -770 -2210
rect -628 -2377 -436 -1815
rect -1388 -2403 -1196 -2402
rect -1024 -2975 -61 -2783
rect -1024 -4497 -832 -2975
rect -253 -4445 -61 -2975
rect -510 -4446 416 -4445
rect -510 -4636 223 -4446
rect 415 -4636 416 -4446
rect -510 -4637 416 -4636
use Comparator  Comparator_0 ../design/JNW_GR05_SKY130A
timestamp 1744491797
transform 1 0 -11 0 1 -5975
box 5350 -4666 13822 1906
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 -72 1 0 2084
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_3
timestamp 1734044400
transform 0 -1 -561 1 0 3382
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_4
timestamp 1734044400
transform 0 -1 728 1 0 2084
box -184 -128 1208 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 -1972 1 0 2084
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1734044400
transform 0 -1 -1972 1 0 784
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1734044400
transform 0 -1 -2772 1 0 784
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1734044400
transform 0 -1 -2772 1 0 2084
box -184 -128 1336 928
use JNWATR_PCH_8C5F0  JNWATR_PCH_8C5F0_1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 -1972 1 0 3384
box -184 -128 1592 928
use JNWATR_PCH_8C5F0  JNWATR_PCH_8C5F0_2
timestamp 1734044400
transform 0 -1 -2772 1 0 3384
box -184 -128 1592 928
use JNWTR_CAPX1  JNWTR_CAPX1_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 -1100 0 1 -5000
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_1
timestamp 1737500400
transform 1 0 -1100 0 1 -3100
box 0 0 1080 1080
use JNWTR_CAPX4  JNWTR_CAPX4_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_TR_SKY130A
timestamp 1744527752
transform 1 0 17728 0 1 -332
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_1
timestamp 1744527752
transform 1 0 4260 0 1 5060
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_2
timestamp 1744527752
transform 1 0 -1580 0 1 -8300
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_3
timestamp 1744527752
transform 1 0 9914 0 1 -170
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_4
timestamp 1744527752
transform 1 0 17004 0 1 -3186
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_5
timestamp 1744527752
transform 1 0 6274 0 1 1536
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_7
timestamp 1744527752
transform 1 0 12484 0 1 -3910
box 480 0 3120 2640
use OTA_Manuel  OTA_Manuel_0 ../design/JNW_GR05_SKY130A
timestamp 1744209957
transform 1 0 -12702 0 1 -4974
box 1600 -402 11980 5848
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1738263620
transform 1 0 -11500 0 1 1000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1738263620
transform 1 0 -11500 0 1 3800
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1738263620
transform 1 0 -10100 0 1 1000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1738263620
transform 1 0 -8700 0 1 1000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1738263620
transform 1 0 -11500 0 1 2400
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1738263620
transform 1 0 -10100 0 1 2400
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1738263620
transform 1 0 -8700 0 1 2400
box 0 0 1340 1340
use JNWATR_NCH_2C1F2  x2 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 2684 0 1 528
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  x4
timestamp 1734044400
transform 0 -1 28 1 0 -4116
box -184 -128 1208 928
use JNWTR_RPPO2  x5 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1743097816
transform 1 0 -7300 0 1 -200
box 0 0 1448 3440
use JNWTR_RPPO16  x10 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1743097816
transform -1 0 -5528 0 -1 7340
box 0 0 4472 3440
<< properties >>
string FIXED_BBOX 0 0 5536 7480
<< end >>
