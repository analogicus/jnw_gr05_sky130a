*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_GR05_lpe.spi
#else
.include ../../../work/xsch/JNW_GR05.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3
.options savecurrents


*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param PERIOD_CLK = 100n
.param vdda = 1.8
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS     VSS      0     dc 0
VDD     VDD_1V8  VSS   dc {vdda}
Vreset  RESET    VSS   dc 0       pulse (0 {vdda} 0  {TRF} {TRF} 50n             590640n      )
VCLK    CLK      VSS   dc 0       pulse (0 {vdda} 0  {TRF} {TRF} {PERIOD_CLK/2}  {PERIOD_CLK} )


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
* .save all
.save i(@m.xdut.x11.x20.xm1.msky130_fd_pr__pfet_01v8[id])

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=14
set color0=white
set color1=black
unset askquit


# write
# -40 -35 -30 -25 -20, -15, -10, -5, 0, 5, 10, 15, 20, 25, 30, 35, 40, 45, 50, 55, 60, 65, 70, 75, 80, 85, 90, 95, 100, 105, 110, 115, 120
set fend = .raw
foreach vtemp -40 
	*-30 -20 -10 0 10 20 30 40 50 60 70 80 90 100 110 120
	option temp=$vtemp
	tran 25n 2.7u 
	write {cicname}_$vtemp$fend
end
quit


.endc

.end
