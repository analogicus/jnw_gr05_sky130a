magic
tech sky130A
magscale 1 2
timestamp 1744469802
<< locali >>
rect 5548 1194 13366 1204
rect 5548 1192 10078 1194
rect 5548 1036 5962 1192
rect 6118 1189 10078 1192
rect 6118 1036 7411 1189
rect 5548 1033 7411 1036
rect 7567 1033 10078 1189
rect 5548 1014 10078 1033
rect 10258 1014 13366 1194
rect 5548 1012 13366 1014
rect 5548 644 5740 1012
rect 6700 628 6892 1012
rect 7008 669 7200 1012
rect 8416 673 8608 1012
rect 9048 666 9240 1012
rect 10456 628 10648 1012
rect 10788 676 10980 1012
rect 11940 676 12132 1012
rect 8289 584 8356 590
rect 8289 529 8295 584
rect 8350 529 8356 584
rect 8289 520 8356 529
rect 8288 468 8356 520
rect 8288 466 8298 468
rect 5548 -358 5740 180
rect 6700 -324 6892 454
rect 9303 328 9370 410
rect 9303 273 9309 328
rect 9364 273 9370 328
rect 9303 267 9370 273
rect 10788 -324 10980 108
rect 11940 -372 12132 220
rect 9311 -481 9369 -475
rect 9311 -527 9317 -481
rect 9363 -527 9369 -481
rect 9311 -638 9369 -527
rect 8283 -738 8339 -685
rect 8283 -782 8289 -738
rect 8333 -782 8339 -738
rect 8283 -788 8339 -782
rect 7388 -1953 7580 -1699
rect 8412 -1953 8604 -1699
rect 9048 -1953 9240 -1700
rect 10072 -1953 10264 -1700
rect 7388 -2008 10265 -1953
rect 7388 -2145 8618 -2008
rect 7388 -2147 7580 -2145
rect 8228 -2384 8420 -2145
rect 8774 -2145 10265 -2008
rect 9252 -2432 9444 -2145
<< viali >>
rect 5962 1036 6118 1192
rect 7411 1033 7567 1189
rect 10078 1014 10258 1194
rect 8295 529 8350 584
rect 9309 273 9364 328
rect 9317 -527 9363 -481
rect 8289 -782 8333 -738
rect 8618 -2164 8774 -2008
<< metal1 >>
rect 5804 1440 13822 1504
rect 5804 674 5868 1440
rect 5956 1192 6124 1204
rect 5956 1036 5962 1192
rect 6118 1036 6124 1192
rect 5956 620 6124 1036
rect 7405 1189 7573 1201
rect 7405 1033 7411 1189
rect 7567 1033 7573 1189
rect 7405 620 7573 1033
rect 10072 1194 10264 1206
rect 10072 1014 10078 1194
rect 10258 1014 10264 1194
rect 8283 584 9562 590
rect 8283 529 8295 584
rect 8350 529 9562 584
rect 8283 523 9562 529
rect 10072 357 10264 1014
rect 11812 686 11876 1440
rect 8095 328 9376 334
rect 8095 273 9309 328
rect 9364 273 9376 328
rect 8095 267 9376 273
rect 5804 -320 5868 123
rect 11812 -290 11876 214
rect 8095 -481 9375 -475
rect 8095 -527 9317 -481
rect 9363 -527 9375 -481
rect 8095 -533 9375 -527
rect 8277 -738 9556 -732
rect 8277 -782 8289 -738
rect 8333 -782 9556 -738
rect 8277 -788 9556 -782
rect 7772 -1320 7964 -874
rect 9304 -948 9368 -942
rect 8284 -960 8348 -954
rect 8284 -1158 8348 -1024
rect 9304 -1156 9368 -1012
rect 9688 -1284 9880 -901
rect 8028 -1842 8220 -1387
rect 8923 -1842 9024 -1841
rect 9432 -1842 9624 -1324
rect 8028 -1943 9624 -1842
rect 8028 -1944 8220 -1943
rect 8612 -2008 8780 -1996
rect 8612 -2164 8618 -2008
rect 8774 -2164 8780 -2008
rect 8612 -2440 8780 -2164
rect 8868 -2464 9060 -1943
rect 9432 -1944 9624 -1943
<< via1 >>
rect 8284 -1024 8348 -960
rect 9304 -1012 9368 -948
<< metal2 >>
rect 9304 1905 9368 1906
rect 7790 1902 8284 1905
rect 7790 1841 8348 1902
rect 8284 -960 8348 1841
rect 9304 1841 9908 1905
rect 9304 -948 9368 1841
rect 8278 -1024 8284 -960
rect 8348 -1024 8354 -960
rect 9298 -1012 9304 -948
rect 9368 -1012 9374 -948
rect 8284 -1154 8348 -1024
use JNWTR_IVX1_CV  x1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1744212116
transform 1 0 5050 0 1 -2180
box -150 -120 2130 440
use JNWTR_IVX1_CV  x2
timestamp 1744212116
transform 1 0 10650 0 1 -2080
box -150 -120 2130 440
use JNWTR_IVX1_CV  x12
timestamp 1744212116
transform 1 0 8150 0 1 -4580
box -150 -120 2130 440
use JNWTR_IVX1_CV  x13
timestamp 1744212116
transform -1 0 9330 0 -1 -3660
box -150 -120 2130 440
use JNWATR_NCH_4C5F0  x14 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1744065478
transform 1 0 10384 0 1 -3272
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  x15
timestamp 1744065478
transform 1 0 5384 0 1 -3272
box -184 -128 1336 928
use JNWTR_CAPX1  x20 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 5300 0 1 -4600
box 0 0 1080 1080
use JNWTR_CAPX1  x21
timestamp 1737500400
transform 1 0 10600 0 1 -4600
box 0 0 1080 1080
use JNWTR_CAPX1  xbuf1
timestamp 1737500400
transform 1 0 7102 0 1 -3273
box 0 0 1080 1080
use JNWTR_CAPX1  xbuf2
timestamp 1737500400
transform 1 0 9600 0 1 -3300
box 0 0 1080 1080
use JNWTR_CAPX1  xbuf3
timestamp 1737500400
transform 1 0 6200 0 1 -1000
box 0 0 1080 1080
use JNWTR_CAPX1  xbuf4
timestamp 1737500400
transform 1 0 10400 0 1 -1000
box 0 0 1080 1080
use JNWATR_NCH_2C1F2  xeval1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 8324 0 1 -3032
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch1
timestamp 1734044400
transform -1 0 8508 0 -1 -1051
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch2
timestamp 1734044400
transform 1 0 9144 0 1 -1852
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch3
timestamp 1734044400
transform 1 0 7484 0 1 -1032
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch4
timestamp 1734044400
transform -1 0 10168 0 -1 -232
box -184 -128 1208 928
use JNWATR_PCH_4C1F2  xpre1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 5644 0 1 -972
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xpre2
timestamp 1734044400
transform 1 0 5644 0 1 28
box -184 -128 1336 928
use JNWATR_PCH_8C1F2  xpre3 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 7104 0 1 28
box -184 -128 1592 928
use JNWATR_PCH_8C1F2  xpre4
timestamp 1734044400
transform -1 0 10552 0 -1 828
box -184 -128 1592 928
use JNWATR_PCH_4C1F2  xpre5
timestamp 1734044400
transform -1 0 12036 0 -1 828
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xpre6
timestamp 1734044400
transform -1 0 12036 0 -1 -172
box -184 -128 1336 928
<< labels >>
flabel metal1 5804 1440 11044 1504 0 FreeSans 1600 0 0 0 CLK
port 6 nsew
flabel metal2 9304 1841 9908 1905 0 FreeSans 1600 0 0 0 Vin2
port 8 nsew
flabel metal2 7790 1841 8284 1905 0 FreeSans 1600 0 0 0 Vin1
port 10 nsew
flabel locali 11358 1012 13366 1204 0 FreeSans 1600 0 0 0 VDD
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 19740 5720
<< end >>
