magic
tech sky130A
magscale 1 2
timestamp 1744466840
<< locali >>
rect 5548 1035 12132 1129
rect 5548 937 6759 1035
rect 5548 655 5740 937
rect 6700 843 6759 937
rect 6939 1029 9474 1035
rect 6939 849 8448 1029
rect 8628 937 9474 1029
rect 8628 849 9239 937
rect 6939 843 9239 849
rect 9654 1029 12132 1035
rect 9654 849 10446 1029
rect 10626 937 11945 1029
rect 10626 849 10980 937
rect 9654 843 10980 849
rect 6700 782 7197 843
rect 8416 816 9239 843
rect 6700 664 7116 782
rect 8416 676 9196 816
rect 10456 676 10980 843
rect 11940 849 11945 937
rect 12125 849 12132 1029
rect 11940 628 12132 849
rect 6724 180 7200 196
rect 5548 -336 5740 180
rect 6700 4 7200 180
rect 8416 116 9048 180
rect 6700 -376 6892 4
rect 8604 -12 9048 116
rect 10456 -12 10980 180
rect 9310 -122 9774 -58
rect 8282 -460 8346 -454
rect 8282 -512 8288 -460
rect 8340 -512 8346 -460
rect 8282 -759 8346 -512
rect 8540 -812 8604 -432
rect 9310 -525 9362 -122
rect 10788 -356 10980 -12
rect 11940 -256 12132 228
rect 5548 -1505 5740 -820
rect 7388 -1285 7580 -879
rect 7686 -1147 8348 -1141
rect 7686 -1199 8290 -1147
rect 8342 -1199 8348 -1147
rect 7686 -1205 8348 -1199
rect 8412 -1337 8604 -842
rect 9048 -1331 9240 -873
rect 9304 -1208 9958 -1144
rect 9304 -1498 9368 -1208
rect 10072 -1285 10264 -832
rect 5548 -1697 7132 -1505
rect 5544 -1910 5659 -1908
rect 5544 -1914 5740 -1910
rect 5544 -1966 5550 -1914
rect 5602 -1966 5740 -1914
rect 5544 -1970 5740 -1966
rect 5544 -1972 5659 -1970
rect 5287 -2046 5480 -1988
rect 6456 -2041 6541 -1697
rect 6940 -1872 7132 -1697
rect 10304 -1596 11216 -1404
rect 11940 -1547 12132 -802
rect 4953 -2408 5145 -2189
rect 5287 -2238 5870 -2046
rect 6196 -2089 6541 -2041
rect 7388 -1984 7580 -1820
rect 10072 -1984 10264 -1820
rect 7388 -1986 10264 -1984
rect 10304 -1986 10496 -1596
rect 11940 -1739 12718 -1547
rect 11245 -1870 11492 -1810
rect 10670 -1950 10980 -1890
rect 11254 -1975 11477 -1930
rect 12042 -1943 12102 -1739
rect 11254 -1986 11310 -1975
rect 11433 -1986 11477 -1975
rect 7388 -1998 11477 -1986
rect 11780 -1989 12102 -1943
rect 6196 -2101 7000 -2089
rect 6196 -2105 6256 -2101
rect 6338 -2105 7000 -2101
rect 6196 -2165 7001 -2105
rect 7388 -2176 11476 -1998
rect 11780 -2013 12600 -1989
rect 11780 -2017 11840 -2013
rect 11957 -2017 12600 -2013
rect 11780 -2040 12600 -2017
rect 11780 -2077 12620 -2040
rect 5287 -2408 5480 -2238
rect 8228 -2385 8420 -2176
rect 4953 -2600 5480 -2408
rect 9252 -2432 9444 -2176
rect 10072 -2178 11476 -2176
rect 12540 -2103 12620 -2077
rect 12640 -2103 12720 -2040
rect 5288 -2672 5480 -2600
rect 6905 -3305 7102 -3097
rect 6903 -3306 7102 -3305
rect 8228 -3306 8420 -2880
rect 9252 -3306 9444 -2848
rect 10288 -3306 10480 -3093
rect 11404 -3130 11596 -3104
rect 11404 -3306 11632 -3130
rect 5287 -3317 9816 -3306
rect 5287 -3497 5678 -3317
rect 5858 -3339 9816 -3317
rect 5858 -3495 8628 -3339
rect 8784 -3495 9816 -3339
rect 5858 -3497 9816 -3495
rect 5287 -3498 9816 -3497
rect 9996 -3309 11404 -3306
rect 9996 -3489 10678 -3309
rect 10858 -3489 11404 -3309
rect 9996 -3498 11404 -3489
rect 11584 -3498 11807 -3306
rect 5287 -3503 9420 -3498
rect 10288 -3503 10480 -3498
rect 6903 -3513 7100 -3503
rect 9240 -3700 9420 -3503
rect 7285 -3940 7429 -3756
rect 7950 -3930 8141 -3870
rect 8201 -3930 8362 -3870
rect 7285 -4004 7440 -3940
rect 7259 -4084 7440 -4004
rect 7285 -4134 7429 -4084
rect 8087 -4121 8205 -3987
rect 8087 -4166 8240 -4121
rect 8060 -4226 8240 -4166
rect 8087 -4300 8240 -4226
rect 8180 -4336 8240 -4300
rect 8420 -4450 8480 -3887
rect 8570 -3930 8782 -3870
rect 8970 -4170 9030 -3790
rect 8618 -4230 9030 -4170
rect 8970 -4361 9030 -4230
rect 12540 -4261 12720 -2103
rect 9226 -4370 9554 -4310
rect 9268 -4484 9518 -4448
rect 10058 -4484 12720 -4261
rect 9268 -4534 12720 -4484
rect 9267 -4605 12720 -4534
rect 9267 -4606 10150 -4605
rect 12540 -4608 12720 -4605
<< viali >>
rect 6759 843 6939 1035
rect 8448 849 8628 1029
rect 9474 843 9654 1035
rect 10446 849 10626 1029
rect 11945 849 12125 1029
rect 9774 -122 9826 -58
rect 8288 -512 8340 -460
rect 9320 -645 9365 -600
rect 7634 -1205 7686 -1141
rect 8290 -1199 8342 -1147
rect 9958 -1208 10010 -1144
rect 5550 -1966 5602 -1914
rect 11216 -1596 11396 -1404
rect 11197 -1870 11245 -1810
rect 6905 -3097 7102 -2912
rect 5678 -3497 5858 -3317
rect 8628 -3495 8784 -3339
rect 9816 -3498 9996 -3306
rect 10678 -3489 10858 -3309
rect 11404 -3498 11584 -3306
rect 6903 -3698 7100 -3513
rect 7902 -3930 7950 -3870
rect 7285 -4266 7429 -4134
rect 8205 -4121 8327 -3987
rect 8782 -3930 8830 -3870
rect 8570 -4230 8618 -4170
rect 9554 -4370 9602 -4310
<< metal1 >>
rect 6753 1035 6945 1047
rect 9468 1035 9660 1047
rect 4606 980 6759 1035
rect 4604 843 6759 980
rect 6939 1029 9474 1035
rect 6939 849 8448 1029
rect 8628 849 9474 1029
rect 6939 843 9474 849
rect 9654 1029 12137 1035
rect 9654 849 10446 1029
rect 10626 849 11945 1029
rect 12125 849 12137 1029
rect 9654 843 12137 849
rect 4604 561 4796 843
rect 4598 369 4604 561
rect 4796 369 4802 561
rect 4917 -1141 4981 -1135
rect 4343 -1205 4917 -1141
rect 4917 -1211 4981 -1205
rect 5804 -1308 5868 234
rect 5932 -700 6124 843
rect 6753 831 6945 843
rect 7392 300 7584 843
rect 9468 831 9660 843
rect 9502 666 9635 718
rect 9687 666 9693 718
rect 6314 26 6506 204
rect 7258 68 7264 132
rect 7328 68 7334 132
rect 8032 26 8224 396
rect 10072 324 10264 843
rect 6314 -166 7722 26
rect 7914 -166 8224 26
rect 9432 196 9624 260
rect 9432 4 9604 196
rect 9432 -4 9624 4
rect 9425 -80 9431 -4
rect 5956 -932 6124 -700
rect 4269 -1372 6019 -1308
rect 6083 -1372 6089 -1308
rect 5801 -1831 5868 -1372
rect 5538 -1914 5614 -1908
rect 5538 -1966 5550 -1914
rect 5602 -1966 5614 -1914
rect 5538 -1972 5614 -1966
rect 5544 -2603 5608 -1972
rect 5801 -2275 5865 -1831
rect 6316 -1985 6508 -212
rect 8032 -556 8224 -166
rect 8282 -144 9431 -80
rect 8282 -460 8346 -144
rect 9425 -196 9431 -144
rect 9623 -196 9629 -4
rect 9768 -58 9832 -46
rect 10328 -58 10392 132
rect 9768 -122 9774 -58
rect 9826 -122 10392 -58
rect 9768 -134 9832 -122
rect 8282 -512 8288 -460
rect 8340 -512 8346 -460
rect 8282 -524 8346 -512
rect 9432 -536 9624 -196
rect 9814 -263 9904 -257
rect 9689 -353 9814 -263
rect 9814 -359 9904 -353
rect 8188 -600 9377 -594
rect 8188 -645 9320 -600
rect 9365 -645 9377 -600
rect 8188 -651 9377 -645
rect 7772 -868 7964 -800
rect 9682 -896 9688 -704
rect 9880 -896 9886 -704
rect 7628 -1141 7692 -1129
rect 6585 -1205 6591 -1141
rect 6655 -1205 7634 -1141
rect 7686 -1205 7692 -1141
rect 7628 -1217 7692 -1205
rect 7772 -1430 7964 -1060
rect 8284 -1147 8348 -1135
rect 8284 -1199 8290 -1147
rect 8342 -1199 8348 -1147
rect 8284 -1276 8348 -1199
rect 9688 -1404 9880 -896
rect 11044 -1018 11108 328
rect 11172 -700 11364 843
rect 11464 718 11516 724
rect 11516 666 11680 718
rect 11464 660 11516 666
rect 11436 -353 11442 -263
rect 11532 -353 11697 -263
rect 11038 -1081 11044 -1018
rect 11107 -1081 11113 -1018
rect 11044 -1085 11108 -1081
rect 9952 -1144 10016 -1132
rect 9952 -1208 9958 -1144
rect 10010 -1204 12756 -1144
rect 10010 -1208 11210 -1204
rect 9952 -1220 10016 -1208
rect 11402 -1208 12756 -1204
rect 11210 -1404 11402 -1396
rect 8028 -1982 8220 -1508
rect 9432 -1982 9624 -1508
rect 11210 -1596 11216 -1404
rect 11396 -1596 11402 -1404
rect 11210 -1608 11402 -1596
rect 11191 -1810 11251 -1798
rect 10555 -1812 11197 -1810
rect 8028 -1985 8612 -1982
rect 6316 -2174 8612 -1985
rect 8804 -2174 9624 -1982
rect 10544 -1870 11197 -1812
rect 11245 -1870 11251 -1810
rect 6316 -2177 8235 -2174
rect 5800 -2339 8548 -2275
rect 8868 -2464 9060 -2174
rect 10544 -2623 10608 -1870
rect 11191 -1882 11251 -1870
rect 6905 -2649 7102 -2643
rect 5672 -3317 5864 -2887
rect 6905 -2906 7102 -2846
rect 6893 -2912 7114 -2906
rect 6893 -3097 6905 -2912
rect 7102 -3097 7114 -2912
rect 6893 -3103 7114 -3097
rect 5672 -3497 5678 -3317
rect 5858 -3497 5864 -3317
rect 5672 -3509 5864 -3497
rect 6112 -3870 6172 -3103
rect 8622 -3279 8790 -2824
rect 7296 -3339 9768 -3279
rect 7296 -3495 8628 -3339
rect 8784 -3495 9768 -3339
rect 6696 -3704 6702 -3507
rect 6899 -3513 7112 -3507
rect 6899 -3698 6903 -3513
rect 7100 -3698 7112 -3513
rect 7296 -3545 9768 -3495
rect 9810 -3306 10002 -3294
rect 9810 -3498 9816 -3306
rect 9996 -3498 10004 -3306
rect 10196 -3498 10202 -3306
rect 10672 -3309 10864 -2956
rect 10672 -3489 10678 -3309
rect 10858 -3489 10864 -3309
rect 9810 -3510 10002 -3498
rect 10672 -3501 10864 -3489
rect 6899 -3704 7112 -3698
rect 8056 -3744 8092 -3741
rect 8013 -3745 8097 -3744
rect 7896 -3870 7956 -3858
rect 6112 -3930 7902 -3870
rect 7950 -3930 7956 -3870
rect 7896 -3942 7956 -3930
rect 8013 -4121 8140 -3745
rect 4598 -4313 4604 -4121
rect 4796 -4134 8140 -4121
rect 8199 -3987 8333 -3545
rect 8524 -3778 8790 -3545
rect 8199 -4121 8205 -3987
rect 8327 -4121 8333 -3987
rect 8199 -4133 8333 -4121
rect 4796 -4266 7285 -4134
rect 7429 -4266 8140 -4134
rect 8564 -4170 8624 -4158
rect 8264 -4230 8270 -4170
rect 8330 -4230 8570 -4170
rect 8618 -4230 8624 -4170
rect 8564 -4242 8624 -4230
rect 4796 -4313 8140 -4266
rect 8702 -4453 8740 -3778
rect 8776 -3870 8836 -3858
rect 8776 -3930 8782 -3870
rect 8830 -3930 9670 -3870
rect 9730 -3930 9736 -3870
rect 8776 -3942 8836 -3930
rect 9548 -4310 9608 -4298
rect 11135 -4310 11195 -3083
rect 11398 -3300 11590 -3294
rect 11392 -3504 11398 -3300
rect 11590 -3504 11596 -3300
rect 11398 -3510 11590 -3504
rect 9548 -4370 9554 -4310
rect 9602 -4370 11195 -4310
rect 9548 -4382 9608 -4370
rect 8702 -4529 8976 -4453
<< via1 >>
rect 4604 369 4796 561
rect 4917 -1205 4981 -1141
rect 9635 666 9687 718
rect 7264 68 7328 132
rect 7722 -166 7914 26
rect 6019 -1372 6083 -1308
rect 9431 -196 9623 -4
rect 9814 -353 9904 -263
rect 7772 -1060 7964 -868
rect 9688 -896 9880 -704
rect 6591 -1205 6655 -1141
rect 11464 666 11516 718
rect 11442 -353 11532 -263
rect 11044 -1081 11107 -1018
rect 11210 -1396 11402 -1204
rect 6905 -2846 7102 -2649
rect 6702 -3704 6899 -3507
rect 10004 -3498 10196 -3306
rect 4604 -4313 4796 -4121
rect 8270 -4230 8330 -4170
rect 9670 -3930 9730 -3870
rect 11398 -3306 11590 -3300
rect 11398 -3498 11404 -3306
rect 11404 -3498 11584 -3306
rect 11584 -3498 11590 -3306
rect 11398 -3504 11590 -3498
<< metal2 >>
rect 9635 718 9687 724
rect 9687 666 11464 718
rect 11516 666 11522 718
rect 9635 660 9687 666
rect 4604 561 4796 567
rect 4604 -4121 4796 369
rect 7264 132 7328 138
rect 7264 62 7328 68
rect 7722 26 7914 32
rect 7470 -166 7479 26
rect 7661 -166 7722 26
rect 9604 2 9796 4
rect 7722 -172 7914 -166
rect 9431 -4 9796 2
rect 9623 -196 10014 -4
rect 10196 -196 10205 -4
rect 9431 -202 9623 -196
rect 11442 -263 11532 -257
rect 9808 -353 9814 -263
rect 9904 -353 11442 -263
rect 11442 -359 11532 -353
rect 9688 -704 9880 -698
rect 7190 -1060 7772 -868
rect 7964 -1060 7970 -868
rect 9880 -896 10214 -704
rect 10396 -896 10405 -704
rect 9688 -902 9880 -896
rect 11210 -1004 11402 -995
rect 11044 -1018 11107 -1012
rect 7190 -1089 7382 -1060
rect 6591 -1141 6655 -1135
rect 4911 -1205 4917 -1141
rect 4981 -1205 6591 -1141
rect 6591 -1211 6655 -1205
rect 7190 -1280 7382 -1271
rect 6019 -1308 6083 -1302
rect 11044 -1308 11107 -1081
rect 11210 -1204 11402 -1186
rect 11038 -1309 11107 -1308
rect 6083 -1372 11107 -1309
rect 6019 -1378 6083 -1372
rect 11204 -1396 11210 -1204
rect 11402 -1396 11408 -1204
rect 6905 -2408 7102 -2399
rect 6905 -2649 7102 -2595
rect 6899 -2846 6905 -2649
rect 7102 -2846 7108 -2649
rect 11398 -3300 11590 -3294
rect 10004 -3306 10196 -3300
rect 10196 -3498 10214 -3306
rect 10396 -3498 10405 -3306
rect 11195 -3498 11204 -3306
rect 11386 -3498 11398 -3306
rect 6702 -3507 6899 -3501
rect 10004 -3504 10196 -3498
rect 6493 -3704 6502 -3507
rect 6689 -3704 6702 -3507
rect 11398 -3510 11590 -3504
rect 6702 -3710 6899 -3704
rect 9670 -3870 9730 -3864
rect 9730 -3930 9874 -3870
rect 9930 -3930 9939 -3870
rect 9670 -3936 9730 -3930
rect 8270 -4170 8330 -4164
rect 6561 -4230 6570 -4170
rect 6626 -4230 8270 -4170
rect 8270 -4236 8330 -4230
rect 4604 -4319 4796 -4313
<< via2 >>
rect 7479 -166 7661 26
rect 10014 -196 10196 -4
rect 10214 -896 10396 -704
rect 7190 -1271 7382 -1089
rect 11210 -1186 11402 -1004
rect 6905 -2595 7102 -2408
rect 10214 -3498 10396 -3306
rect 11204 -3498 11386 -3306
rect 6502 -3704 6689 -3507
rect 9874 -3930 9930 -3870
rect 6570 -4230 6626 -4170
<< metal3 >>
rect 7474 26 7666 31
rect 7051 -166 7479 26
rect 7661 -166 7666 26
rect 7474 -171 7666 -166
rect 10009 -4 10201 1
rect 10009 -196 10014 -4
rect 10196 -196 10596 -4
rect 10009 -201 10201 -196
rect 10209 -704 10401 -699
rect 10209 -896 10214 -704
rect 10396 -896 10401 -704
rect 7185 -1089 7387 -1084
rect 6905 -1264 7102 -1258
rect 7185 -1271 7190 -1089
rect 7382 -1271 7387 -1089
rect 7185 -1276 7387 -1271
rect 6905 -2193 7102 -1459
rect 7190 -1496 7382 -1276
rect 7190 -1692 7382 -1686
rect 10209 -1906 10401 -896
rect 11210 -999 11402 -604
rect 11205 -1004 11407 -999
rect 11205 -1186 11210 -1004
rect 11402 -1186 11407 -1004
rect 11205 -1191 11407 -1186
rect 10209 -2102 10401 -2096
rect 6905 -2403 7488 -2193
rect 6900 -2408 7488 -2403
rect 6900 -2595 6905 -2408
rect 7102 -2595 7107 -2408
rect 6900 -2600 7107 -2595
rect 10209 -3306 10401 -3004
rect 10209 -3498 10214 -3306
rect 10396 -3498 10401 -3306
rect 6497 -3506 6694 -3502
rect 10209 -3503 10401 -3498
rect 11199 -3306 11391 -3301
rect 11199 -3498 11204 -3306
rect 11386 -3498 11391 -3306
rect 6202 -3507 6694 -3506
rect 6202 -3703 6502 -3507
rect 6497 -3704 6502 -3703
rect 6689 -3704 6694 -3507
rect 6497 -3709 6694 -3704
rect 11199 -3796 11391 -3498
rect 9869 -3870 9935 -3865
rect 10162 -3870 10168 -3868
rect 9869 -3930 9874 -3870
rect 9930 -3930 10168 -3870
rect 9869 -3935 9935 -3930
rect 10162 -3932 10168 -3930
rect 10232 -3932 10238 -3868
rect 6362 -4232 6368 -4168
rect 6432 -4170 6438 -4168
rect 6565 -4170 6631 -4165
rect 6432 -4230 6570 -4170
rect 6626 -4230 6631 -4170
rect 6432 -4232 6438 -4230
rect 6565 -4235 6631 -4230
<< via3 >>
rect 6905 -1459 7102 -1264
rect 7190 -1686 7382 -1496
rect 10209 -2096 10401 -1906
rect 10168 -3932 10232 -3868
rect 6368 -4232 6432 -4168
<< metal4 >>
rect 6905 -1263 7102 -681
rect 6904 -1264 7103 -1263
rect 6904 -1459 6905 -1264
rect 7102 -1459 7103 -1264
rect 6904 -1460 7103 -1459
rect 7189 -1496 7383 -1495
rect 7189 -1686 7190 -1496
rect 7382 -1686 7383 -1496
rect 7189 -1687 7383 -1686
rect 7190 -2366 7382 -1687
rect 10208 -1906 10402 -1905
rect 10208 -2096 10209 -1906
rect 10401 -2096 10402 -1906
rect 10208 -2097 10402 -2096
rect 10209 -2596 10401 -2097
rect 10167 -3868 10233 -3867
rect 10167 -3932 10168 -3868
rect 10232 -3870 10233 -3868
rect 10232 -3930 12230 -3870
rect 10232 -3932 10233 -3930
rect 10167 -3933 10233 -3932
rect 6367 -4168 6433 -4167
rect 6367 -4170 6368 -4168
rect 6070 -4230 6368 -4170
rect 6367 -4232 6368 -4230
rect 6432 -4232 6433 -4168
rect 6367 -4233 6433 -4232
rect 12170 -4530 12230 -3930
use JNWTR_IVX1_CV  x1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1744212116
transform 1 0 5050 0 1 -2180
box -150 -120 2130 440
use JNWTR_IVX1_CV  x2
timestamp 1744212116
transform 1 0 10650 0 1 -2080
box -150 -120 2130 440
use JNWTR_IVX1_CV  x12
timestamp 1744212116
transform 1 0 8150 0 1 -4580
box -150 -120 2130 440
use JNWTR_IVX1_CV  x13
timestamp 1744212116
transform -1 0 9330 0 -1 -3660
box -150 -120 2130 440
use JNWATR_NCH_4C5F0  x14 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1744065478
transform 1 0 10384 0 1 -3272
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  x15
timestamp 1744065478
transform 1 0 5384 0 1 -3272
box -184 -128 1336 928
use JNWTR_CAPX1  x20 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 5300 0 1 -4600
box 0 0 1080 1080
use JNWTR_CAPX1  x21
timestamp 1737500400
transform 1 0 10600 0 1 -4600
box 0 0 1080 1080
use JNWTR_CAPX1  xbuf1
timestamp 1737500400
transform 1 0 7102 0 1 -3273
box 0 0 1080 1080
use JNWTR_CAPX1  xbuf2
timestamp 1737500400
transform 1 0 9600 0 1 -3300
box 0 0 1080 1080
use JNWTR_CAPX1  xbuf3
timestamp 1737500400
transform 1 0 6200 0 1 -1000
box 0 0 1080 1080
use JNWTR_CAPX1  xbuf4
timestamp 1737500400
transform 1 0 10400 0 1 -1000
box 0 0 1080 1080
use JNWATR_NCH_2C1F2  xeval1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 8324 0 1 -3032
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch1
timestamp 1734044400
transform -1 0 8508 0 -1 -1172
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch2
timestamp 1734044400
transform 1 0 9144 0 1 -1972
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch3
timestamp 1734044400
transform 1 0 7484 0 1 -1032
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch4
timestamp 1734044400
transform -1 0 10168 0 -1 -232
box -184 -128 1208 928
use JNWATR_PCH_4C1F2  xpre1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 5644 0 1 -972
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xpre2
timestamp 1734044400
transform 1 0 5644 0 1 28
box -184 -128 1336 928
use JNWATR_PCH_8C1F2  xpre3 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 7104 0 1 28
box -184 -128 1592 928
use JNWATR_PCH_8C1F2  xpre4
timestamp 1734044400
transform -1 0 10552 0 -1 828
box -184 -128 1592 928
use JNWATR_PCH_4C1F2  xpre5
timestamp 1734044400
transform 1 0 10884 0 1 28
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xpre6
timestamp 1734044400
transform 1 0 10884 0 1 -972
box -184 -128 1336 928
<< labels >>
flabel metal1 10010 -1208 10596 -1144 0 FreeSans 1600 0 0 0 Vin2
port 0 nsew
flabel metal1 6948 -1205 7634 -1141 0 FreeSans 1600 0 0 0 Vin1
port 2 nsew
flabel locali 5288 -3498 11404 -3306 0 FreeSans 1600 0 0 0 VSS
port 10 nsew
flabel metal1 4751 -1372 4843 -1308 0 FreeSans 1600 0 0 0 CLK
port 4 nsew
flabel metal4 12170 -4530 12230 -3870 0 FreeSans 1600 0 0 0 Vout
port 12 nsew
flabel metal1 4843 843 11364 1035 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 19740 5720
<< end >>
