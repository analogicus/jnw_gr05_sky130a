magic
tech sky130A
magscale 1 2
timestamp 1744209957
<< locali >>
rect 11788 5433 11980 5438
rect 4598 5292 11980 5433
rect 4562 4743 4719 5008<
rect 7434 4706 11032 4898
rect 4562 4087 4719 4093
rect 4562 3942 4568 4087
rect 4713 3942 4719 4087
rect 4912 4072 5024 4544
rect 4562 3665 4719 3942
rect 5488 403 5680 1580
rect 6206 446 7088 452
rect 6206 394 7030 446
rect 7082 394 7088 446
rect 6206 388 7088 394
rect 7152 361 7344 1584
rect 4572 143 4708 352
rect 5488 -204 5680 -20
rect 5488 -374 6774 -204
rect 7152 -204 7344 9
rect 7520 -204 7712 4706
rect 10840 4562 11032 4706
rect 8564 3796 9018 3802
rect 8564 3712 8928 3796
rect 9012 3712 9018 3796
rect 8564 3706 9018 3712
rect 11788 3616 11980 5292
rect 7888 3608 11980 3616
rect 7888 3428 8278 3608
rect 8458 3606 11980 3608
rect 8458 3428 10078 3606
rect 7888 3426 10078 3428
rect 10258 3426 11980 3606
rect 7888 3424 11980 3426
rect 7888 3236 8080 3424
rect 8202 3196 8674 3230
rect 7888 1928 8068 2694
rect 9040 2020 9232 2828
rect 9688 1951 9880 2729
rect 10840 1982 11032 2828
rect 9040 1206 9232 1506
rect 9690 1240 9882 1474
rect 9690 1234 10264 1240
rect 9690 1054 10078 1234
rect 10258 1054 10264 1234
rect 9690 1048 10264 1054
rect 7888 -204 8080 180
rect 9040 -204 9232 183
rect 9688 -204 9880 180
rect 10840 -100 11032 180
rect 10840 -204 11034 -100
rect 6954 -207 11034 -204
rect 6954 -374 8668 -207
rect 5488 -375 8668 -374
rect 8836 -208 11034 -207
rect 8836 -375 10078 -208
rect 5488 -388 10078 -375
rect 10258 -388 11034 -208
rect 5488 -396 11034 -388
rect 5488 -402 5680 -396
<< viali >>
rect 4562 4598 4719 4743
rect 4568 3942 4713 4087
rect 6154 388 6206 452
rect 7030 394 7082 446
rect 4572 19 4708 143
rect 6774 -374 6954 -194
rect 8480 3706 8564 3802
rect 8928 3712 9012 3796
rect 8278 3428 8458 3608
rect 10078 3426 10258 3606
rect 8150 3196 8202 3230
rect 8674 3196 8708 3230
rect 9040 1026 9232 1206
rect 10078 1054 10258 1234
rect 8668 -375 8836 -207
rect 10078 -388 10258 -208
<< metal1 >>
rect 7326 5032 8208 5096
rect 4550 4743 4731 4749
rect 4550 4598 4562 4743
rect 4719 4598 4731 4743
rect 8144 4624 8208 5032
rect 9944 5036 10926 5100
rect 9944 4607 10008 5036
rect 4550 4592 4731 4598
rect 4562 4087 4719 4592
rect 4562 3942 4568 4087
rect 4713 3942 4719 4087
rect 4562 3930 4719 3942
rect 8323 3811 8436 4076
rect 5842 3802 8436 3811
rect 8474 3802 8570 3814
rect 5842 3706 8480 3802
rect 8564 3706 8570 3802
rect 5842 3698 8436 3706
rect 5872 1872 6064 3698
rect 8474 3694 8570 3706
rect 8272 3608 8464 3620
rect 8272 3428 8278 3608
rect 8458 3428 8464 3608
rect 8144 2336 8208 2808
rect 8272 2740 8464 3428
rect 8656 3230 8848 4208
rect 10118 3802 10214 4066
rect 8916 3796 10214 3802
rect 8916 3712 8928 3796
rect 9012 3712 10214 3796
rect 8916 3706 10214 3712
rect 8656 3196 8674 3230
rect 8708 3196 8848 3230
rect 8656 3150 8848 3196
rect 10072 3606 10264 3618
rect 10072 3426 10078 3606
rect 10258 3426 10264 3606
rect 10072 2968 10264 3426
rect 10456 3116 10648 4196
rect 9944 2578 10008 2762
rect 10492 2578 10556 2836
rect 9944 2514 10556 2578
rect 8316 2336 8976 2340
rect 8144 2276 8976 2336
rect 8144 2272 8380 2276
rect 8912 1904 8976 2276
rect 9944 2034 10008 2514
rect 6148 452 6212 464
rect 6768 452 6960 1814
rect 7024 524 7088 1728
rect 8272 934 8464 1560
rect 8656 1218 8848 1632
rect 10072 1234 10264 1640
rect 8656 1212 9224 1218
rect 8656 1206 9244 1212
rect 8656 1026 9040 1206
rect 9232 1026 9244 1206
rect 10072 1054 10078 1234
rect 10258 1054 10264 1234
rect 10072 1042 10264 1054
rect 10456 1182 10648 1618
rect 9028 1020 9244 1026
rect 10456 990 11584 1182
rect 8272 870 8976 934
rect 8272 604 8464 870
rect 8912 732 8976 870
rect 8912 724 10008 732
rect 8916 668 10008 724
rect 10456 568 10648 990
rect 5874 388 6154 452
rect 6206 388 6212 452
rect 6148 376 6212 388
rect 7024 446 7088 486
rect 7024 394 7030 446
rect 7082 394 7088 446
rect 4560 143 4720 149
rect 4560 19 4572 143
rect 4708 105 4720 143
rect 4708 19 6017 105
rect 4560 13 6017 19
rect 4561 7 6017 13
rect 6768 -194 6960 380
rect 7024 372 7088 394
rect 6768 -374 6774 -194
rect 6954 -374 6960 -194
rect 6768 -386 6960 -374
rect 8662 -207 8842 395
rect 8912 211 10008 275
rect 10072 -202 10264 332
rect 8662 -375 8668 -207
rect 8836 -375 8842 -207
rect 8662 -387 8842 -375
rect 10066 -208 10270 -202
rect 10066 -388 10078 -208
rect 10258 -388 10270 -208
rect 10066 -394 10270 -388
use JNWTR_RPPO2  x5 ../JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1743097816
transform 0 1 1600 -1 0 5848
box 0 0 1448 3440
use JNWTR_RPPO16  x6 ../JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1743097816
transform 0 1 1600 -1 0 4272
box 0 0 4472 3440
use JNWATR_PCH_12C5F0  xb1 ../JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1744194304
transform -1 0 7248 0 -1 628
box -184 -128 1848 928
use JNWATR_PCH_12C5F0  xb2
timestamp 1744194304
transform -1 0 7248 0 -1 2228
box -184 -128 1848 928
use JNWATR_NCH_4C5F0  xli1 ../JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1744065478
transform 1 0 7984 0 1 2628
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xli2 ../JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 7984 0 1 3928
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xlo1
timestamp 1744065478
transform -1 0 9136 0 -1 2128
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xlo2 ../JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform -1 0 9136 0 -1 828
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xri1
timestamp 1744065478
transform 1 0 9784 0 1 2628
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xri2
timestamp 1734044400
transform 1 0 9784 0 1 3928
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xro1
timestamp 1744065478
transform 1 0 9784 0 1 1328
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xro2
timestamp 1734044400
transform 1 0 9784 0 1 28
box -184 -128 1336 928
<< labels >>
flabel metal1 7326 5032 8208 5096 0 FreeSans 1600 0 0 0 V_n
port 2 nsew
flabel metal1 9944 5036 10926 5100 0 FreeSans 1600 0 0 0 V_p
port 3 nsew
flabel locali 11788 3424 11980 5438 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
flabel metal1 10456 990 11584 1182 0 FreeSans 1600 0 0 0 I_out
port 9 nsew
flabel locali 10258 -396 11034 -204 0 FreeSans 1600 0 0 0 VDD
port 15 nsew
<< properties >>
string FIXED_BBOX 0 0 8944 5640
<< end >>
