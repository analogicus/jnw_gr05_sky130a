magic
tech sky130A
magscale 1 2
timestamp 1744572521
<< locali >>
rect -10229 7451 -2855 7452
rect -10229 7187 1768 7451
rect -10229 6190 -9964 7187
rect -10229 5747 -9964 5937
rect -10229 5057 -9964 5494
rect -11437 4902 -9964 5057
rect -5585 6821 1768 7187
rect -5585 6568 1086 6821
rect 1339 6568 1768 6821
rect -5585 6104 1768 6568
rect -5585 5912 2594 6104
rect -5585 5528 2358 5912
rect -5585 5275 1091 5528
rect 1344 5458 2358 5528
rect 1344 5278 2140 5458
rect 2320 5278 2358 5458
rect 1344 5275 2358 5278
rect -5585 5080 2358 5275
rect -5585 4954 2628 5080
rect -11437 4066 -11282 4902
rect -10387 4066 -10232 4902
rect -11437 4061 -10232 4066
rect -10229 4104 -9964 4902
rect -5628 4888 2628 4954
rect -5628 4831 1768 4888
rect -5628 4696 -3387 4831
rect -9563 4180 -9396 4420
rect -6172 4180 -5991 4420
rect -5628 4104 -3697 4696
rect -10229 4061 -3697 4104
rect -11437 4027 -3697 4061
rect -3081 4310 1768 4831
rect -3081 4027 -1583 4310
rect -11437 3989 -1583 4027
rect -11437 3928 -10232 3989
rect -10229 3928 -1583 3989
rect -11473 3920 -1583 3928
rect -11473 3887 -6464 3920
rect -11475 3839 -6464 3887
rect -11475 3637 -8051 3839
rect -11469 3459 -8051 3637
rect -7872 3667 -6464 3839
rect -6211 3667 -1583 3920
rect -7872 3480 -1583 3667
rect -525 4212 1768 4310
rect -525 3480 1005 4212
rect -7872 3459 1005 3480
rect -11469 2646 -11280 3459
rect -10416 3330 -10061 3459
rect -10416 3008 -10040 3330
rect -10421 2646 -10040 3008
rect -9985 2686 -9846 3459
rect -8990 3388 -8487 3459
rect -8990 2690 -8851 3388
rect -9985 2646 -9839 2686
rect -9021 2646 -8851 2690
rect -8815 2661 -8487 3388
rect -7614 3140 1005 3459
rect -7614 2673 -7425 3140
rect -8815 2646 -8439 2661
rect -7621 2646 -7425 2673
rect -7420 2646 -7279 3140
rect -6896 2942 -6444 2948
rect -6896 2762 -6890 2942
rect -6710 2762 -6444 2942
rect -6896 2756 -6444 2762
rect -11469 2627 -7279 2646
rect -11405 2458 -7279 2627
rect -11473 2108 -7279 2458
rect -11473 2079 -7754 2108
rect -11474 1303 -11262 2031
rect -10421 1876 -9839 2031
rect -11474 1257 -11239 1303
rect -10421 1261 -9876 1876
rect -9021 1445 -8439 2079
rect -7621 1782 -7425 2108
rect -9021 1261 -8474 1445
rect -10421 1260 -8243 1261
rect -7614 1260 -7425 1782
rect -10421 1257 -7425 1260
rect -11474 1183 -7425 1257
rect -11474 1125 -7465 1183
rect -7420 1125 -7279 2108
rect -5884 1848 -4513 3140
rect -1465 3012 1005 3140
rect 1561 3325 2090 3371
rect 1561 3145 1678 3325
rect 1858 3145 2090 3325
rect 1561 3041 2090 3145
rect -1465 2180 -915 3012
rect 1561 2180 1891 3041
rect -11474 1071 -7279 1125
rect -11474 1068 -9937 1071
rect -11474 1058 -11239 1068
rect -11474 1027 -11162 1058
rect -10285 1027 -9937 1068
rect -9015 1027 -7279 1071
rect -11474 858 -7279 1027
rect -11476 823 -7279 858
rect -11476 792 -7268 823
rect -11476 746 -10942 792
rect -11474 -461 -10982 746
rect -7773 -51 -7268 792
rect -5882 752 -4513 1848
rect -2172 1840 -741 2180
rect -413 2174 2050 2180
rect -413 1940 751 2174
rect -413 1840 538 1940
rect 745 1846 751 1940
rect 1079 1846 2050 2174
rect 3211 2146 3403 3370
rect 745 1840 2050 1846
rect -3612 752 -3420 880
rect -5882 737 -2930 752
rect -2463 737 -2172 752
rect -5882 688 -2172 737
rect -1466 688 538 1840
rect 1561 832 1891 1840
rect -5882 396 538 688
rect 1005 826 1891 832
rect 1005 646 1011 826
rect 1191 646 1891 826
rect 1005 640 1891 646
rect -5882 318 -5741 396
rect -5630 380 538 396
rect -5630 362 -2930 380
rect -4764 318 -2930 362
rect -2463 318 538 380
rect -7773 -268 -5895 -51
rect -5393 -76 -5193 -72
rect -4281 -76 -4089 -6
rect -1466 34 538 318
rect -5550 -243 -5076 -76
rect -7773 -444 -7408 -268
rect -7790 -461 -7408 -444
rect -11474 -770 -7408 -461
rect -11474 -4974 -10982 -770
rect -7773 -902 -7408 -770
rect -11480 -5106 -10982 -4974
rect -7717 -5106 -7408 -902
rect -5550 -2258 -4990 -243
rect -1466 -374 -16 34
rect 392 -374 538 34
rect -1466 -852 538 -374
rect -1466 -1032 -628 -852
rect -436 -1032 538 -852
rect -1466 -1250 538 -1032
rect -1466 -1358 -22 -1250
rect -2058 -1550 -22 -1358
rect -7214 -2580 -4990 -2258
rect -1759 -1658 -22 -1550
rect 398 -1658 538 -1250
rect -1759 -2233 538 -1658
rect 1561 -2055 1891 640
rect 7938 -1572 9228 -1152
rect -1759 -2513 58 -2233
rect -7214 -2901 -7022 -2580
rect -5550 -2999 -4990 -2580
rect -1670 -2641 58 -2513
rect 466 -2527 538 -2233
rect 1560 -2418 1962 -2055
rect 1560 -2428 2052 -2418
rect 466 -2641 539 -2527
rect -1670 -2693 539 -2641
rect -1862 -2719 539 -2693
rect -1862 -2978 -1670 -2719
rect 1560 -2920 6588 -2428
rect -1754 -2996 -1734 -2978
rect -11480 -5178 -7408 -5106
rect -7214 -5220 -7022 -5178
rect -5546 -5220 -4993 -2999
rect -1810 -3188 -1734 -2996
rect -664 -3188 -604 -3060
rect -172 -3188 543 -3060
rect -1862 -3642 -1734 -3494
rect 351 -3636 543 -3188
rect -129 -3642 543 -3636
rect -1862 -3686 -845 -3642
rect -1111 -3822 -845 -3686
rect -129 -3822 -123 -3642
rect 57 -3670 543 -3642
rect 57 -3822 223 -3670
rect -1111 -4020 -667 -3822
rect -129 -3828 223 -3822
rect 100 -3850 223 -3828
rect 415 -3850 543 -3670
rect 100 -4020 543 -3850
rect -1111 -4212 543 -4020
rect 1560 -5220 2052 -2920
rect 8808 -3477 9228 -1572
rect 7504 -3897 9228 -3477
rect -7214 -5584 2052 -5220
<< viali >>
rect -10229 5937 -9964 6190
rect -10229 5494 -9964 5747
rect 1086 6568 1339 6821
rect 1091 5275 1344 5528
rect 2140 5278 2320 5458
rect -9791 4180 -9563 4420
rect -5991 4180 -5763 4420
rect -6464 3667 -6211 3920
rect -6890 2762 -6710 2942
rect -6444 2756 -6264 2948
rect 1678 3145 1858 3325
rect -741 1840 -413 2180
rect 751 1846 1079 2174
rect 1011 646 1191 826
rect -4281 -6 -4089 174
rect -16 -374 392 34
rect -628 -1032 -436 -852
rect -22 -1658 398 -1250
rect -1862 -2693 -1670 -2513
rect 58 -2641 466 -2233
rect -845 -3822 -665 -3642
rect -123 -3822 57 -3642
rect 223 -3850 415 -3670
rect 7096 -3897 7504 -3477
<< metal1 >>
rect 712 6827 977 6833
rect 977 6821 1351 6827
rect 977 6568 1086 6821
rect 1339 6568 1351 6821
rect 977 6562 1351 6568
rect 712 6556 977 6562
rect -10228 6521 -9963 6527
rect -10228 6196 -9963 6256
rect -10241 6190 -9952 6196
rect -10241 5937 -10229 6190
rect -9964 5937 -9952 6190
rect -10241 5931 -9952 5937
rect 1162 5887 1354 5893
rect -10241 5747 -9952 5753
rect -10241 5494 -10229 5747
rect -9964 5494 -9952 5747
rect -10241 5488 -9952 5494
rect 687 5534 952 5540
rect 1162 5534 1354 5695
rect -10228 5443 -9963 5488
rect 952 5528 1356 5534
rect 2107 5528 2113 5720
rect 2305 5528 2660 5720
rect 952 5275 1091 5528
rect 1344 5275 1356 5528
rect 952 5269 1356 5275
rect 2128 5458 2956 5464
rect 2128 5278 2140 5458
rect 2320 5278 2956 5458
rect 2128 5272 2956 5278
rect 687 5263 952 5269
rect -10228 5172 -9963 5178
rect -5994 4909 -5787 4915
rect -5994 4504 -5787 4702
rect 1162 4684 1354 5269
rect 9184 5208 9190 5267
rect 2955 5144 9190 5208
rect 9184 5075 9190 5144
rect 9382 5075 9388 5267
rect -9797 4420 -9557 4432
rect -10984 4180 -9791 4420
rect -9563 4180 -9557 4420
rect -6001 4420 -2564 4504
rect 1162 4454 1354 4492
rect 3766 4454 3830 4460
rect -6001 4312 -5991 4420
rect -9797 4168 -9557 4180
rect -5997 4180 -5991 4312
rect -5763 4312 -2564 4420
rect -2228 4390 3766 4454
rect -5763 4180 -4516 4312
rect -5997 4168 -5757 4180
rect 1162 4118 1354 4390
rect 3766 4384 3830 4390
rect -6051 3926 -5786 3932
rect -1185 3926 1402 4118
rect 1594 4071 1600 4118
rect 3777 4071 3841 4077
rect 1594 4007 3777 4071
rect 1594 3926 1600 4007
rect 3777 4001 3841 4007
rect -6476 3920 -6051 3926
rect -6476 3667 -6464 3920
rect -6211 3667 -6051 3920
rect -6476 3661 -6051 3667
rect -3397 3672 -2434 3864
rect -2311 3862 -960 3864
rect -2311 3672 -1929 3862
rect -1935 3670 -1929 3672
rect -1737 3672 -960 3862
rect -1737 3670 -1731 3672
rect -6051 3655 -5786 3661
rect -3387 3606 -1535 3608
rect -3387 3544 -1164 3606
rect -1599 3542 -1164 3544
rect -1599 3444 -1535 3542
rect -1604 3381 -1535 3444
rect -10859 2900 -9478 3092
rect -6450 2948 -6258 2960
rect -10859 1648 -10667 2900
rect -9670 1648 -9478 2900
rect -7896 2942 -6444 2948
rect -7896 2762 -6890 2942
rect -6710 2762 -6444 2942
rect -7896 2756 -6444 2762
rect -6264 2756 -3304 2948
rect -3096 2756 -2404 2948
rect -6450 2744 -6258 2756
rect -4558 1863 -4494 2756
rect -1604 2564 -1540 3381
rect 1311 3331 1503 3337
rect 1503 3325 1870 3331
rect 1503 3145 1678 3325
rect 1858 3145 1870 3325
rect 1503 3139 1870 3145
rect 1311 3133 1503 3139
rect 1480 2820 1672 2844
rect -418 2628 264 2820
rect 398 2628 1672 2820
rect -3110 2372 -1929 2564
rect -1737 2372 -492 2564
rect -446 2372 388 2564
rect -1604 2308 -1540 2372
rect 1480 2308 1672 2628
rect -2932 2244 -768 2308
rect -202 2244 126 2308
rect 553 2244 1672 2308
rect -4564 1799 -4558 1863
rect -4494 1799 -4488 1863
rect -10859 1456 -3260 1648
rect -2999 1456 -2540 1648
rect -4558 1245 -4494 1251
rect -4558 58 -4494 1181
rect -4281 832 -4089 838
rect -4281 180 -4089 640
rect -4293 174 -4077 180
rect -4293 -6 -4281 174
rect -4089 -6 -4077 174
rect -3900 114 -3836 1456
rect -2304 1261 -1740 1264
rect -2304 1072 -1929 1261
rect -1935 1069 -1929 1072
rect -1737 1069 -1731 1261
rect -1604 1008 -1540 2244
rect -747 2180 -407 2192
rect -747 1840 -741 2180
rect -413 2174 1091 2180
rect -413 1846 751 2174
rect 1079 1846 1091 2174
rect -413 1840 1091 1846
rect -747 1828 -407 1840
rect -3042 944 -1532 1008
rect 643 832 835 838
rect -3414 557 -3284 749
rect 835 826 1203 832
rect 835 646 1011 826
rect 1191 646 1203 826
rect 835 640 1203 646
rect 643 634 835 640
rect -3900 62 -2758 114
rect -3900 50 -2694 62
rect -4293 -12 -4077 -6
rect -22 34 398 46
rect -22 -374 -16 34
rect 392 -374 398 34
rect -22 -539 398 -374
rect -640 -852 -424 -846
rect -640 -1032 -628 -852
rect -436 -1032 -424 -852
rect -640 -1038 -424 -1032
rect -628 -1133 -436 -1038
rect -22 -1244 398 -959
rect -628 -1331 -436 -1325
rect -34 -1250 410 -1244
rect -34 -1658 -22 -1250
rect 398 -1658 410 -1250
rect -34 -1664 410 -1658
rect -1862 -2210 -1670 -2204
rect 575 -2227 995 -2221
rect -1862 -2507 -1670 -2402
rect 46 -2233 575 -2227
rect -1874 -2513 -1658 -2507
rect -1874 -2693 -1862 -2513
rect -1670 -2693 -1658 -2513
rect 46 -2641 58 -2233
rect 466 -2641 575 -2233
rect 46 -2647 575 -2641
rect 575 -2653 995 -2647
rect -1874 -2699 -1658 -2693
rect -664 -3380 -478 -3374
rect 1480 -3380 1672 2244
rect 8900 -1028 9190 -836
rect 9382 -1028 9388 -836
rect -664 -3572 -478 -3566
rect -318 -3572 1672 -3380
rect 7090 -3477 7510 -3465
rect -857 -3642 69 -3636
rect -857 -3822 -845 -3642
rect -665 -3822 -123 -3642
rect 57 -3822 69 -3642
rect -857 -3828 69 -3822
rect 211 -3670 427 -3664
rect 211 -3850 223 -3670
rect 415 -3850 427 -3670
rect 211 -3856 427 -3850
rect -1282 -3956 -550 -3892
rect 223 -3909 415 -3856
rect 5354 -3897 5360 -3477
rect 5780 -3897 7096 -3477
rect 7504 -3897 7510 -3477
rect 7090 -3909 7510 -3897
rect 223 -4107 415 -4101
<< via1 >>
rect 712 6562 977 6827
rect -10228 6256 -9963 6521
rect 1162 5695 1354 5887
rect -10228 5178 -9963 5443
rect 687 5269 952 5534
rect 2113 5528 2305 5720
rect -5994 4702 -5787 4909
rect 9190 5075 9382 5267
rect 1162 4492 1354 4684
rect 3766 4390 3830 4454
rect 1402 3926 1594 4118
rect 3777 4007 3841 4071
rect -6051 3661 -5786 3926
rect -1929 3670 -1737 3862
rect 1311 3139 1503 3331
rect -1929 2372 -1737 2564
rect -4558 1799 -4494 1863
rect -4558 1181 -4494 1245
rect -4281 640 -4089 832
rect -1929 1069 -1737 1261
rect 643 640 835 832
rect -22 -959 398 -539
rect -628 -1325 -436 -1133
rect -1862 -2402 -1670 -2210
rect 575 -2647 995 -2227
rect 9190 -1028 9382 -836
rect -664 -3566 -478 -3380
rect 5360 -3897 5780 -3477
rect 223 -4101 415 -3909
<< metal2 >>
rect -10228 6822 -9963 6831
rect 304 6827 559 6831
rect -10228 6521 -9963 6567
rect 299 6822 712 6827
rect 299 6567 304 6822
rect 559 6567 712 6822
rect 299 6562 712 6567
rect 977 6562 983 6827
rect 304 6558 559 6562
rect -10234 6256 -10228 6521
rect -9963 6256 -9957 6521
rect 1162 6229 1354 6238
rect 1162 5887 1354 6047
rect 1156 5695 1162 5887
rect 1354 5695 1360 5887
rect 2113 5720 2305 5726
rect 340 5534 595 5538
rect 335 5529 687 5534
rect -10234 5178 -10228 5443
rect -9963 5178 -9957 5443
rect 335 5274 340 5529
rect 595 5274 687 5529
rect 335 5269 687 5274
rect 952 5269 958 5534
rect 1793 5528 1802 5720
rect 1984 5528 2113 5720
rect 2113 5522 2305 5528
rect 340 5265 595 5269
rect 9190 5267 9382 5273
rect -5994 5179 -5787 5188
rect -10228 5153 -9963 5178
rect -5994 4909 -5787 4982
rect 1142 5052 1374 5061
rect -10228 4889 -9963 4898
rect -6000 4702 -5994 4909
rect -5787 4702 -5781 4909
rect 1142 4684 1374 4830
rect 1142 4492 1162 4684
rect 1354 4492 1374 4684
rect 1142 4472 1374 4492
rect 1402 4434 1594 4443
rect 3760 4390 3766 4454
rect 3830 4390 5718 4454
rect 1402 4118 1594 4252
rect -5673 3926 -5418 3930
rect 3771 4007 3777 4071
rect 3841 4007 4204 4071
rect 5654 3994 5718 4390
rect -6057 3661 -6051 3926
rect -5786 3921 -5412 3926
rect -5786 3666 -5673 3921
rect -5418 3666 -5412 3921
rect 1402 3920 1594 3926
rect -5786 3661 -5412 3666
rect -1929 3862 -1737 3868
rect -5673 3657 -5418 3661
rect -1929 3331 -1737 3670
rect -1929 3139 1311 3331
rect 1503 3139 1509 3331
rect -1929 2564 -1737 3139
rect -4558 1863 -4494 1869
rect -4558 1245 -4494 1799
rect -1929 1261 -1737 2372
rect -4564 1181 -4558 1245
rect -4494 1181 -4488 1245
rect -1929 832 -1737 1069
rect -4287 640 -4281 832
rect -4089 640 643 832
rect 835 640 841 832
rect -28 -959 -22 -539
rect 398 -959 1508 -539
rect -634 -1325 -628 -1133
rect -436 -1325 -430 -1133
rect -628 -1388 -436 -1325
rect -628 -1579 -436 -1570
rect -1868 -2402 -1862 -2210
rect -1670 -2402 -1583 -2210
rect -1401 -2402 -1392 -2210
rect 1088 -2227 1508 -959
rect 9190 -836 9382 5075
rect 9190 -1034 9382 -1028
rect 569 -2647 575 -2227
rect 995 -2647 1508 -2227
rect -1014 -3572 -1005 -3380
rect -823 -3566 -664 -3380
rect -478 -3566 -262 -3380
rect -86 -3566 -77 -3380
rect 1088 -3477 1508 -2647
rect 5360 -3477 5780 -3471
rect -823 -3572 -637 -3566
rect 1088 -3897 5360 -3477
rect 5360 -3903 5780 -3897
rect 217 -4101 223 -3909
rect 415 -4101 421 -3909
rect 223 -4151 415 -4101
rect 223 -4342 415 -4333
<< via2 >>
rect -10228 6567 -9963 6822
rect 304 6567 559 6822
rect 1162 6047 1354 6229
rect 340 5274 595 5529
rect 1802 5528 1984 5720
rect -10228 4898 -9963 5153
rect -5994 4982 -5787 5179
rect 1142 4830 1374 5052
rect 1402 4252 1594 4434
rect -5673 3666 -5418 3921
rect -628 -1570 -436 -1388
rect -1583 -2402 -1401 -2210
rect -1005 -3572 -823 -3380
rect -262 -3566 -86 -3380
rect 223 -4333 415 -4151
<< metal3 >>
rect -3402 6827 -3137 6968
rect -1937 6827 -1672 6953
rect -10233 6822 564 6827
rect -10233 6567 -10228 6822
rect -9963 6567 304 6822
rect 559 6567 564 6822
rect -10233 6562 564 6567
rect 1162 6645 1354 6651
rect -9405 6536 -7720 6562
rect -9405 5158 -9140 6536
rect -7985 5158 -7720 6536
rect -4836 5534 -4571 6562
rect -3402 5534 -3137 6562
rect -1937 5534 -1672 6562
rect -441 5534 -176 6562
rect 1162 6234 1354 6455
rect 1157 6229 1359 6234
rect 1157 6047 1162 6229
rect 1354 6047 1359 6229
rect 1157 6042 1359 6047
rect 1797 5720 1989 5725
rect -4836 5529 600 5534
rect -4836 5274 340 5529
rect 595 5274 600 5529
rect 1512 5528 1518 5720
rect 1708 5528 1802 5720
rect 1984 5528 1989 5720
rect 1797 5523 1989 5528
rect -4836 5269 600 5274
rect 1142 5470 1374 5476
rect -10233 5153 -7720 5158
rect -10233 4898 -10228 5153
rect -9963 4898 -7720 5153
rect -6566 4977 -6560 5184
rect -6355 5179 -5782 5184
rect -6355 4982 -5994 5179
rect -5787 4982 -5782 5179
rect -6355 4977 -5782 4982
rect -10233 4893 -7720 4898
rect -4836 4268 -4571 5269
rect -3402 4268 -3137 5269
rect -1937 4268 -1672 5269
rect -452 4268 -176 5269
rect 1142 5057 1374 5240
rect 1137 5052 1379 5057
rect 1137 4830 1142 5052
rect 1374 4830 1379 5052
rect 1137 4825 1379 4830
rect -4953 4003 -176 4268
rect 1397 4434 1599 4439
rect 1397 4252 1402 4434
rect 1594 4252 1599 4434
rect 1397 4247 1599 4252
rect -4953 3926 -4571 4003
rect -5678 3921 -4571 3926
rect -5678 3666 -5673 3921
rect -5418 3666 -4571 3921
rect -5678 3661 -4571 3666
rect -4836 2859 -4571 3661
rect -3402 2941 -3137 4003
rect -1937 2941 -1672 4003
rect -3402 2859 -1672 2941
rect -441 2859 -176 4003
rect 1402 3906 1594 4247
rect 1402 3710 1594 3716
rect -4836 2594 -176 2859
rect -633 -1388 -431 -1383
rect -633 -1570 -628 -1388
rect -436 -1570 -431 -1388
rect -633 -1575 -431 -1570
rect -628 -1624 -436 -1575
rect -628 -1820 -436 -1814
rect -1588 -2210 -1396 -2205
rect -1588 -2402 -1583 -2210
rect -1401 -2402 -1387 -2210
rect -1197 -2402 -1191 -2210
rect -1588 -2407 -1396 -2402
rect -1010 -3380 -818 -2752
rect -1010 -3572 -1005 -3380
rect -823 -3572 -818 -3380
rect -1010 -4017 -818 -3572
rect -267 -3380 -81 -2782
rect -267 -3566 -262 -3380
rect -86 -3566 -81 -3380
rect -267 -4089 -81 -3566
rect 218 -4151 420 -4146
rect 218 -4333 223 -4151
rect 415 -4333 420 -4151
rect 218 -4338 420 -4333
rect 223 -4446 415 -4338
rect 223 -4642 415 -4636
<< via3 >>
rect 1162 6455 1354 6645
rect 1518 5528 1708 5720
rect -6560 4977 -6355 5184
rect 1142 5240 1374 5470
rect 1402 3716 1594 3906
rect -628 -1814 -436 -1624
rect -1387 -2402 -1197 -2210
rect 223 -4636 415 -4446
<< metal4 >>
rect -1984 6978 -209 7065
rect -4962 6786 -209 6978
rect -9426 6514 -7595 6721
rect -9426 5093 -9219 6514
rect -7802 5184 -7595 6514
rect -6561 5184 -6354 5185
rect -7802 5093 -6560 5184
rect -9426 4977 -6560 5093
rect -6355 4977 -6353 5184
rect -9426 4886 -7489 4977
rect -6561 4976 -6354 4977
rect -4962 4807 -4770 6786
rect -3302 5415 -3110 6786
rect -1984 5415 -1792 6786
rect -426 6646 -209 6786
rect -426 6645 1355 6646
rect -426 6455 1162 6645
rect 1354 6633 1355 6645
rect 1354 6455 1709 6633
rect -426 6454 1709 6455
rect -426 5471 -209 6454
rect -28 6441 1709 6454
rect 1517 5720 1709 6441
rect 1517 5528 1518 5720
rect 1708 5528 1709 5720
rect 1517 5499 1709 5528
rect 67 5471 1709 5499
rect -452 5470 1709 5471
rect -452 5415 1142 5470
rect -4738 5240 1142 5415
rect 1374 5307 1709 5470
rect 1374 5240 1375 5307
rect -4738 5239 1375 5240
rect -4738 5223 -209 5239
rect -4738 4807 -4546 5223
rect -4962 4615 -4546 4807
rect -4962 3907 -4770 4615
rect -4738 3907 -4546 4615
rect -3302 3907 -3110 5223
rect -1984 3907 -1792 5223
rect -401 3907 -209 5223
rect 1517 3907 1709 5307
rect -4962 3906 1709 3907
rect -4962 3716 1402 3906
rect 1594 3716 1709 3906
rect -4962 3715 1709 3716
rect -4738 2667 -4546 3715
rect -3302 2667 -3110 3715
rect -1984 2667 -1792 3715
rect -401 2667 -209 3715
rect 9 3709 1709 3715
rect -4738 2475 -209 2667
rect -3302 2469 -1792 2475
rect -629 -1624 -435 -1623
rect -629 -1814 -628 -1624
rect -436 -1814 -435 -1624
rect -629 -1815 -435 -1814
rect -1388 -2210 -1196 -2209
rect -1388 -2402 -1387 -2210
rect -1197 -2402 -770 -2210
rect -628 -2377 -436 -1815
rect -1388 -2403 -1196 -2402
rect -1024 -2975 -61 -2783
rect -1024 -4497 -832 -2975
rect -253 -4445 -61 -2975
rect -510 -4446 416 -4445
rect -510 -4636 223 -4446
rect 415 -4636 416 -4446
rect -510 -4637 416 -4636
use Comparator  Comparator_0 ../design/JNW_GR05_SKY130A
timestamp 1744491797
transform 1 0 -3650 0 1 2166
box 5350 -4666 13822 1906
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 -72 1 0 2084
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_3
timestamp 1734044400
transform 0 -1 -561 1 0 3382
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_4
timestamp 1734044400
transform 0 -1 728 1 0 2084
box -184 -128 1208 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 -1972 1 0 2084
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1734044400
transform 0 -1 -1972 1 0 784
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1734044400
transform 0 -1 -2772 1 0 784
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1734044400
transform 0 -1 -2772 1 0 2084
box -184 -128 1336 928
use JNWATR_PCH_8C5F0  JNWATR_PCH_8C5F0_1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 -1972 1 0 3384
box -184 -128 1592 928
use JNWATR_PCH_8C5F0  JNWATR_PCH_8C5F0_2
timestamp 1734044400
transform 0 -1 -2772 1 0 3384
box -184 -128 1592 928
use JNWTR_CAPX1  JNWTR_CAPX1_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 -1100 0 1 -5000
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_1
timestamp 1737500400
transform 1 0 -1100 0 1 -3100
box 0 0 1080 1080
use JNWTR_CAPX4  JNWTR_CAPX4_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_TR_SKY130A
timestamp 1744527752
transform 1 0 -2880 0 1 4800
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_1
timestamp 1744527752
transform 1 0 -5780 0 1 -800
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_2
timestamp 1744527752
transform 1 0 -2880 0 1 2000
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_3
timestamp 1744527752
transform 1 0 -5780 0 1 4800
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_4
timestamp 1744527752
transform 1 0 -10280 0 1 4500
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_6
timestamp 1744527752
transform 1 0 -2880 0 1 -800
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_7
timestamp 1744527752
transform 1 0 -5780 0 1 2000
box 480 0 3120 2640
use OTA_Manuel  OTA_Manuel_0 ../design/JNW_GR05_SKY130A
timestamp 1744209957
transform 1 0 -12702 0 1 -4974
box 1600 -402 11980 5848
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1738263620
transform 1 0 -11500 0 1 1000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1738263620
transform 1 0 -11500 0 1 3800
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1738263620
transform 1 0 -10100 0 1 1000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1738263620
transform 1 0 -8700 0 1 1000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1738263620
transform 1 0 -11500 0 1 2400
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1738263620
transform 1 0 -10100 0 1 2400
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1738263620
transform 1 0 -8700 0 1 2400
box 0 0 1340 1340
use JNWATR_NCH_2C1F2  x2 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 3228 1 0 4984
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  x4
timestamp 1734044400
transform 0 -1 28 1 0 -4116
box -184 -128 1208 928
use JNWTR_RPPO2  x5 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1743097816
transform 1 0 -7300 0 1 -200
box 0 0 1448 3440
use JNWTR_RPPO16  x10 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1743097816
transform -1 0 -5528 0 -1 7340
box 0 0 4472 3440
<< labels >>
flabel locali -3081 4310 1768 7451 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel space -3866 -5370 -2624 -5178 0 FreeSans 1600 0 0 0 VDD_1V8
port 3 nsew
flabel space 4898 3606 10172 3670 0 FreeSans 1600 0 0 0 CLK
port 5 nsew
flabel space 7406 -1028 9286 -836 0 FreeSans 1600 0 0 0 CompOut
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 5536 7480
<< end >>
