magic
tech sky130A
magscale 1 2
timestamp 1744533318
<< locali >>
rect -2139 3140 771 3332
rect -6896 2942 -6444 2948
rect -6896 2762 -6890 2942
rect -6710 2762 -6444 2942
rect -6896 2756 -6444 2762
rect -11474 1092 -11375 2525
rect -10421 2151 -10349 2696
rect -9911 2525 -9839 2686
rect -9021 2525 -8949 2690
rect -10320 2426 -8535 2525
rect -10074 2248 -9975 2426
rect -9911 2151 -9839 2426
rect -9021 2151 -8949 2426
rect -8674 2229 -8575 2426
rect -8511 2151 -8439 2661
rect -10421 2079 -7754 2151
rect -10421 1261 -10349 2079
rect -9911 1876 -9839 2079
rect -9021 1261 -8949 2079
rect -8511 1445 -8439 2079
rect -7621 1782 -7549 2673
rect -2172 1940 773 2180
rect -10421 1189 -8243 1261
rect -10285 1026 -9937 1125
rect -9015 1026 -7386 1125
rect -3612 737 -3420 880
rect -2155 737 968 880
rect -3612 688 968 737
rect -3612 380 -1905 688
rect -856 -2996 -670 -2994
rect -1810 -3188 -670 -2996
rect -664 -3188 -604 -2996
rect -1681 -3494 -670 -3188
rect -1862 -3598 -670 -3494
rect -1862 -3642 -667 -3598
rect -1862 -3686 -845 -3642
rect -1111 -3822 -845 -3686
rect -1111 -4020 -667 -3822
rect -1111 -4212 68 -4020
<< viali >>
rect -6890 2762 -6710 2942
rect -6444 2756 -6264 2948
rect -845 -3822 -665 -3642
<< metal1 >>
rect -10859 2900 -9478 3092
rect -6450 2948 -6258 2960
rect -10859 1648 -10667 2900
rect -9670 1648 -9478 2900
rect -7896 2942 -6444 2948
rect -7896 2762 -6890 2942
rect -6710 2762 -6444 2942
rect -7896 2756 -6444 2762
rect -6264 2756 -3304 2948
rect -3096 2756 -2404 2948
rect -6450 2744 -6258 2756
rect -4558 1863 -4494 2756
rect 398 2628 1672 2820
rect -3096 2372 -2404 2564
rect -434 2372 255 2564
rect -2932 2244 -2468 2308
rect -2132 2244 -768 2308
rect -202 2244 126 2308
rect -4564 1799 -4558 1863
rect -4494 1799 -4488 1863
rect -10859 1456 -3260 1648
rect -2999 1456 -2540 1648
rect -4558 1245 -4494 1251
rect -4558 58 -4494 1181
rect -3900 114 -3836 1456
rect -3112 1072 -2552 1264
rect -1532 1008 -1468 2244
rect -3042 944 -1468 1008
rect -3900 62 -2758 114
rect -3900 50 -2694 62
rect 1480 -3380 1672 2628
rect -318 -3572 1672 -3380
rect -857 -3642 -296 -3636
rect -857 -3822 -845 -3642
rect -665 -3822 -296 -3642
rect -857 -3828 -296 -3822
rect -1282 -3956 -850 -3892
rect -670 -3956 -590 -3892
<< via1 >>
rect -4558 1799 -4494 1863
rect -4558 1181 -4494 1245
<< metal2 >>
rect -4558 1863 -4494 1869
rect -4558 1245 -4494 1799
rect -4564 1181 -4558 1245
rect -4494 1181 -4488 1245
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -5862 0 1 8356
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_1
timestamp 1734044400
transform 0 -1 -72 1 0 2084
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_3
timestamp 1734044400
transform 1 0 -2270 0 1 9144
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_4
timestamp 1734044400
transform 0 -1 728 1 0 2084
box -184 -128 1208 928
use JNWATR_PCH_4C5F0__0  JNWATR_PCH_4C5F0__0_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 -2772 1 0 2084
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  JNWATR_PCH_4C5F0__0_1
timestamp 1734044400
transform 0 -1 -1972 1 0 784
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  JNWATR_PCH_4C5F0__0_2
timestamp 1734044400
transform 0 -1 -2772 1 0 784
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  JNWATR_PCH_4C5F0__0_3
timestamp 1734044400
transform 0 -1 -1972 1 0 2084
box -184 -128 1336 928
use JNWATR_PCH_8C5F0  JNWATR_PCH_8C5F0_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -2992 0 1 7272
box -184 -128 1592 928
use JNWATR_PCH_8C5F0  JNWATR_PCH_8C5F0_1
timestamp 1734044400
transform 1 0 716 0 1 7938
box -184 -128 1592 928
use JNWTR_CAPX1  JNWTR_CAPX1_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 -150 0 1 10082
box 0 0 1080 1080
use JNWTR_CAPX4  JNWTR_CAPX4_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_TR_SKY130A
timestamp 1744527752
transform 1 0 17728 0 1 -332
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_1
timestamp 1744527752
transform 1 0 4260 0 1 5060
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_2
timestamp 1744527752
transform 1 0 -234 0 1 -7799
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_3
timestamp 1744527752
transform 1 0 9914 0 1 -170
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_4
timestamp 1744527752
transform 1 0 17004 0 1 -3186
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_5
timestamp 1744527752
transform 1 0 6274 0 1 1536
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_7
timestamp 1744527752
transform 1 0 12484 0 1 -3910
box 480 0 3120 2640
use JNWTR_RPPO16  JNWTR_RPPO16_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1743097816
transform 1 0 -13900 0 1 7100
box 0 0 4472 3440
use JNWTR_RPPO16  JNWTR_RPPO16_2
timestamp 1743097816
transform 1 0 13172 0 1 5630
box 0 0 4472 3440
use JNWTR_RPPO16  JNWTR_RPPO16_4
timestamp 1743097816
transform 1 0 -6500 0 1 12000
box 0 0 4472 3440
use OTA_Manuel  OTA_Manuel_0 ../design/JNW_GR05_SKY130A
timestamp 1744209957
transform 1 0 -12702 0 1 -4974
box 1600 -402 11980 5848
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1738263620
transform 1 0 -11500 0 1 1000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1738263620
transform 1 0 -9400 0 1 4300
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1738263620
transform 1 0 -10100 0 1 1000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1738263620
transform 1 0 -8700 0 1 1000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1738263620
transform 1 0 -11500 0 1 2400
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1738263620
transform 1 0 -10100 0 1 2400
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1738263620
transform 1 0 -8700 0 1 2400
box 0 0 1340 1340
use JNWATR_NCH_2C1F2  x2 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 3108 0 1 16
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  x4
timestamp 1734044400
transform 0 -1 28 1 0 -4116
box -184 -128 1208 928
use JNWTR_RPPO2  x5 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1743097816
transform 1 0 -7300 0 1 -200
box 0 0 1448 3440
use JNWTR_RPPO8  x7 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1744527752
transform 1 0 -150 0 1 11382
box 0 0 2744 3440
use JNWTR_RPPO16  x10
timestamp 1743097816
transform 1 0 -12900 0 1 12100
box 0 0 4472 3440
<< properties >>
string FIXED_BBOX 0 0 5536 7480
<< end >>
