magic
tech sky130A
magscale 1 2
timestamp 1744491797
<< locali >>
rect 5410 1205 5606 1206
rect 5410 1204 5740 1205
rect 5410 1198 13366 1204
rect 5410 1194 11562 1198
rect 5410 1192 10078 1194
rect 5410 1036 5962 1192
rect 6118 1189 10078 1192
rect 6118 1036 7411 1189
rect 5410 1033 7411 1036
rect 7567 1033 10078 1189
rect 5410 1014 10078 1033
rect 10258 1018 11562 1194
rect 11742 1018 13366 1198
rect 10258 1014 13366 1018
rect 5410 1012 13366 1014
rect 5410 628 5740 1012
rect 6700 628 6892 1012
rect 7008 669 7200 1012
rect 8416 673 8608 1012
rect 9048 666 9240 1012
rect 10456 628 10648 1012
rect 10788 676 10980 1012
rect 11940 676 12132 1012
rect 5410 180 5606 628
rect 8289 584 8356 590
rect 8289 529 8295 584
rect 8350 529 8356 584
rect 8289 520 8356 529
rect 8288 468 8356 520
rect 8288 466 8298 468
rect 5410 -358 5740 180
rect 6700 -324 6892 454
rect 9303 328 9370 410
rect 9303 273 9309 328
rect 9364 273 9370 328
rect 9303 267 9370 273
rect 5410 -545 5606 -358
rect 5410 -1774 5612 -545
rect 5410 -1809 6160 -1774
rect 5410 -4482 5612 -1809
rect 7090 -1892 7210 -164
rect 10788 -324 10980 108
rect 11940 -372 12132 220
rect 9311 -481 9369 -475
rect 9311 -527 9317 -481
rect 9363 -527 9369 -481
rect 9311 -638 9369 -527
rect 8283 -738 8339 -685
rect 8283 -782 8289 -738
rect 8333 -782 8339 -738
rect 8283 -788 8339 -782
rect 11040 -796 11100 -790
rect 11040 -844 11046 -796
rect 11094 -844 11100 -796
rect 7150 -1914 7210 -1892
rect 7388 -1699 7452 -1434
rect 7516 -1699 7580 -1512
rect 7388 -1953 7580 -1699
rect 8412 -1953 8604 -1699
rect 9048 -1953 9240 -1700
rect 10072 -1720 10264 -1700
rect 10072 -1800 10640 -1720
rect 10072 -1848 10620 -1800
rect 10072 -1952 10674 -1848
rect 11040 -1940 11100 -844
rect 11940 -1166 12132 -820
rect 11940 -1358 12724 -1166
rect 12540 -1800 12720 -1358
rect 11670 -1852 11690 -1840
rect 11636 -1854 11700 -1852
rect 10072 -1953 10740 -1952
rect 7388 -1980 10740 -1953
rect 7388 -2008 9868 -1980
rect 7388 -2126 8618 -2008
rect 6138 -2136 8618 -2126
rect 6138 -2316 6528 -2136
rect 6708 -2145 8618 -2136
rect 6708 -2158 8420 -2145
rect 6708 -2258 7893 -2158
rect 8005 -2258 8420 -2158
rect 8774 -2033 9868 -2008
rect 9933 -1991 10740 -1980
rect 9933 -2030 11310 -1991
rect 9933 -2033 10740 -2030
rect 8774 -2145 10740 -2033
rect 6708 -2316 8420 -2258
rect 6138 -2318 8420 -2316
rect 6138 -2368 6330 -2318
rect 8294 -2388 8420 -2318
rect 6138 -2480 6330 -2448
rect 8294 -2500 8334 -2388
rect 9252 -2432 9444 -2145
rect 8294 -2756 8320 -2500
rect 10288 -2624 10480 -2145
rect 11628 -2226 11700 -1854
rect 11820 -2046 12600 -1986
rect 11312 -2290 11700 -2226
rect 11312 -2772 11376 -2290
rect 8294 -2956 8420 -2880
rect 7290 -3000 8420 -2956
rect 7290 -3104 7501 -3000
rect 7593 -3096 8420 -3000
rect 9252 -3083 9444 -2832
rect 9252 -3096 9309 -3083
rect 7593 -3102 9309 -3096
rect 7593 -3104 8618 -3102
rect 7290 -3148 8618 -3104
rect 8156 -3282 8618 -3148
rect 8798 -3151 9309 -3102
rect 9389 -3096 9444 -3083
rect 10416 -3096 10480 -2934
rect 9389 -3151 10480 -3096
rect 8798 -3206 10480 -3151
rect 8798 -3274 8874 -3206
rect 8942 -3274 10480 -3206
rect 8798 -3282 10480 -3274
rect 8156 -3288 10480 -3282
rect 7936 -3350 8708 -3324
rect 7893 -3380 8708 -3350
rect 7936 -3384 8708 -3380
rect 9076 -3361 9256 -3288
rect 9914 -3318 10480 -3288
rect 11440 -3318 11632 -3116
rect 9076 -3393 9106 -3361
rect 9226 -3399 9256 -3361
rect 9896 -3324 12878 -3318
rect 8558 -3510 8618 -3508
rect 8526 -3570 8808 -3510
rect 7816 -4482 7996 -3580
rect 8100 -3940 8180 -3762
rect 8558 -4090 8618 -3570
rect 9436 -3950 9496 -3430
rect 9896 -3504 10678 -3324
rect 10858 -3504 12878 -3324
rect 9896 -3510 12878 -3504
rect 11480 -3736 11625 -3510
rect 9436 -4008 9576 -3950
rect 9458 -4010 9576 -4008
rect 9344 -4482 9509 -4116
rect 10058 -4190 10138 -4180
rect 10058 -4482 10238 -4190
rect 5410 -4621 10238 -4482
rect 5414 -4660 10238 -4621
rect 5414 -4662 10140 -4660
rect 5888 -4666 6252 -4662
<< viali >>
rect 5962 1036 6118 1192
rect 7411 1033 7567 1189
rect 10078 1014 10258 1194
rect 11562 1018 11742 1198
rect 8295 529 8350 584
rect 9309 273 9364 328
rect 7090 -164 7210 -56
rect 9317 -527 9363 -481
rect 8289 -782 8333 -738
rect 11046 -844 11094 -796
rect 6400 -1996 6452 -1944
rect 6528 -2316 6708 -2136
rect 7893 -2258 8005 -2158
rect 8618 -2164 8774 -2008
rect 9868 -2033 9933 -1980
rect 7501 -3104 7593 -3000
rect 8618 -3282 8798 -3102
rect 9309 -3151 9389 -3083
rect 8874 -3274 8942 -3206
rect 8478 -3570 8526 -3510
rect 8100 -3762 8180 -3694
rect 10678 -3504 10858 -3324
rect 11480 -3869 11625 -3736
rect 9576 -4010 9624 -3950
<< metal1 >>
rect 5804 1440 8484 1504
rect 8548 1440 13822 1504
rect 5804 674 5868 1440
rect 5956 1192 6124 1204
rect 5956 1036 5962 1192
rect 6118 1036 6124 1192
rect 5956 620 6124 1036
rect 7405 1189 7573 1201
rect 7405 1033 7411 1189
rect 7567 1033 7573 1189
rect 7405 620 7573 1033
rect 10072 1194 10264 1206
rect 10072 1014 10078 1194
rect 10258 1014 10264 1194
rect 8283 584 9562 590
rect 5804 -320 5868 123
rect 5932 -430 6124 556
rect 8283 529 8295 584
rect 8350 529 9562 584
rect 8283 523 9562 529
rect 6316 24 6508 394
rect 10072 364 10264 1014
rect 11556 1198 11748 1210
rect 11556 1018 11562 1198
rect 11742 1018 11748 1198
rect 8032 334 8224 336
rect 8032 267 8096 334
rect 8163 328 9376 334
rect 8163 273 9309 328
rect 9364 273 9376 328
rect 11556 300 11748 1018
rect 11812 686 11876 1440
rect 8163 267 9376 273
rect 8032 24 8224 267
rect 6316 -56 8224 24
rect 6316 -164 7090 -56
rect 7210 -164 8224 -56
rect 6316 -178 8224 -164
rect 8032 -475 8224 -178
rect 9432 22 9624 260
rect 11172 22 11364 260
rect 9432 -39 11364 22
rect 9432 -117 10094 -39
rect 10172 -117 11364 -39
rect 9432 -178 11364 -117
rect 9432 -406 9624 -178
rect 8032 -481 9375 -475
rect 8032 -482 9317 -481
rect 8095 -527 9317 -482
rect 9363 -527 9375 -481
rect 8095 -533 9375 -527
rect 6316 -1050 6508 -706
rect 8277 -738 9556 -732
rect 8277 -782 8289 -738
rect 8333 -782 9556 -738
rect 8277 -788 9556 -782
rect 11040 -796 11100 -178
rect 11556 -682 11748 178
rect 11812 -290 11876 214
rect 11040 -844 11046 -796
rect 11094 -844 11100 -796
rect 11040 -856 11100 -844
rect 7772 -1050 7964 -874
rect 9304 -948 9368 -942
rect 6316 -1242 7964 -1050
rect 8284 -960 8348 -954
rect 8284 -1158 8348 -1024
rect 9304 -1156 9368 -1012
rect 9688 -1054 9880 -901
rect 11172 -1054 11364 -740
rect 6925 -1401 7052 -1242
rect 7772 -1320 7964 -1242
rect 9688 -1246 11364 -1054
rect 9688 -1284 9880 -1246
rect 6919 -1528 6925 -1401
rect 7052 -1528 7058 -1401
rect 6522 -1860 6858 -1756
rect 8028 -1842 8220 -1387
rect 8923 -1842 9024 -1841
rect 9432 -1842 9624 -1324
rect 10686 -1382 10816 -1376
rect 6394 -1944 6458 -1932
rect 6394 -1996 6400 -1944
rect 6452 -1996 6458 -1944
rect 6394 -2450 6458 -1996
rect 6522 -2136 6714 -1860
rect 8028 -1943 9624 -1842
rect 8028 -1944 8220 -1943
rect 6522 -2316 6528 -2136
rect 6708 -2316 6714 -2136
rect 7893 -1976 8005 -1970
rect 7893 -2152 8005 -2088
rect 8612 -2008 8780 -1996
rect 7881 -2158 8017 -2152
rect 7881 -2258 7893 -2158
rect 8005 -2258 8017 -2158
rect 8612 -2164 8618 -2008
rect 8774 -2164 8780 -2008
rect 7881 -2264 8017 -2258
rect 8484 -2202 8548 -2196
rect 6522 -2670 6714 -2316
rect 8484 -2410 8548 -2266
rect 8612 -2440 8780 -2164
rect 8868 -2464 9060 -1943
rect 9432 -1944 9624 -1943
rect 9868 -1891 9933 -1885
rect 9868 -1974 9933 -1956
rect 9856 -1980 9945 -1974
rect 9856 -2033 9868 -1980
rect 9933 -2033 9945 -1980
rect 9856 -2039 9945 -2033
rect 6927 -3080 7078 -2916
rect 7495 -3000 7599 -2988
rect 7495 -3104 7501 -3000
rect 7593 -3104 7631 -3000
rect 7735 -3104 7741 -3000
rect 8612 -3102 8804 -2568
rect 9309 -2964 9389 -2958
rect 9309 -3077 9389 -3044
rect 7495 -3116 7599 -3104
rect 6927 -3237 7078 -3231
rect 6962 -3501 7029 -3237
rect 8612 -3282 8618 -3102
rect 8798 -3282 8804 -3102
rect 9297 -3083 9401 -3077
rect 9297 -3151 9309 -3083
rect 9389 -3151 9401 -3083
rect 9297 -3157 9401 -3151
rect 8612 -3294 8804 -3282
rect 8868 -3206 8948 -3194
rect 8868 -3274 8874 -3206
rect 8942 -3274 8948 -3206
rect 8472 -3501 8532 -3498
rect 6962 -3510 8532 -3501
rect 6962 -3570 8478 -3510
rect 8526 -3570 8532 -3510
rect 6962 -3577 8532 -3570
rect 8472 -3582 8532 -3577
rect 8868 -3688 8948 -3274
rect 10672 -3324 10864 -2952
rect 11056 -3194 12936 -3002
rect 11102 -3196 11202 -3194
rect 11102 -3302 11202 -3296
rect 10672 -3504 10678 -3324
rect 10858 -3504 10864 -3324
rect 10672 -3516 10864 -3504
rect 8088 -3694 8948 -3688
rect 8088 -3762 8100 -3694
rect 8180 -3762 8948 -3694
rect 8088 -3768 8948 -3762
rect 8868 -4164 8948 -3768
rect 9570 -3950 9630 -3938
rect 11124 -3950 11184 -3302
rect 11217 -3875 11223 -3730
rect 11368 -3736 11637 -3730
rect 11368 -3869 11480 -3736
rect 11625 -3869 11637 -3736
rect 11368 -3875 11637 -3869
rect 9570 -4010 9576 -3950
rect 9624 -4010 11184 -3950
rect 9570 -4022 9630 -4010
<< via1 >>
rect 8484 1440 8548 1504
rect 8096 267 8163 334
rect 10094 -117 10172 -39
rect 8284 -1024 8348 -960
rect 9304 -1012 9368 -948
rect 6925 -1528 7052 -1401
rect 10686 -1376 10816 -1246
rect 7893 -2088 8005 -1976
rect 8484 -2266 8548 -2202
rect 9868 -1956 9933 -1891
rect 6927 -3231 7078 -3080
rect 7631 -3104 7735 -3000
rect 9309 -3044 9389 -2964
rect 11102 -3296 11202 -3196
rect 11223 -3875 11368 -3730
<< metal2 >>
rect 9304 1905 9368 1906
rect 7790 1902 8284 1905
rect 7790 1841 8348 1902
rect 8096 334 8163 340
rect 8096 170 8163 267
rect 8096 104 8163 113
rect 8284 -960 8348 1841
rect 9304 1841 9908 1905
rect 8484 1504 8548 1510
rect 8278 -1024 8284 -960
rect 8348 -1024 8354 -960
rect 8284 -1154 8348 -1024
rect 6925 -1401 7052 -1395
rect 6925 -1593 7052 -1528
rect 6921 -1710 6930 -1593
rect 7047 -1710 7056 -1593
rect 7893 -1615 8005 -1606
rect 6925 -1714 7052 -1710
rect 7893 -1976 8005 -1717
rect 7887 -2088 7893 -1976
rect 8005 -2088 8011 -1976
rect 8484 -2202 8548 1440
rect 9304 -948 9368 1841
rect 10094 -39 10172 -33
rect 9900 -117 9909 -39
rect 9977 -117 10094 -39
rect 10094 -123 10172 -117
rect 9298 -1012 9304 -948
rect 9368 -1012 9374 -948
rect 10680 -1376 10686 -1246
rect 10816 -1376 10822 -1246
rect 10686 -1475 10816 -1376
rect 10686 -1604 10816 -1595
rect 9868 -1677 9933 -1668
rect 9868 -1891 9933 -1733
rect 9862 -1956 9868 -1891
rect 9933 -1956 9939 -1891
rect 8478 -2266 8484 -2202
rect 8548 -2266 8554 -2202
rect 9309 -2846 9389 -2837
rect 9309 -2964 9389 -2916
rect 7631 -3000 7735 -2994
rect 6921 -3231 6927 -3080
rect 7078 -3231 7084 -3080
rect 7735 -3104 7788 -3000
rect 7882 -3104 7891 -3000
rect 9303 -3044 9309 -2964
rect 9389 -3044 9395 -2964
rect 7631 -3110 7735 -3104
rect 6927 -3296 7078 -3231
rect 11096 -3296 11102 -3196
rect 11202 -3296 11208 -3196
rect 11102 -3336 11202 -3296
rect 11102 -3435 11202 -3426
rect 6927 -3446 7078 -3437
rect 11223 -3730 11368 -3724
rect 11000 -3875 11009 -3730
rect 11144 -3875 11223 -3730
rect 11223 -3881 11368 -3875
<< via2 >>
rect 8096 113 8163 170
rect 6930 -1710 7047 -1593
rect 7893 -1717 8005 -1615
rect 9909 -117 9977 -39
rect 10686 -1595 10816 -1475
rect 9868 -1733 9933 -1677
rect 9309 -2916 9389 -2846
rect 7788 -3104 7882 -3000
rect 6927 -3437 7078 -3296
rect 11102 -3426 11202 -3336
rect 11009 -3875 11144 -3730
<< metal3 >>
rect 8091 170 8168 175
rect 8091 113 8096 170
rect 8163 113 8168 170
rect 8091 108 8168 113
rect 8096 43 8163 108
rect 8096 -28 8163 -22
rect 9904 -39 9982 -34
rect 9780 -117 9786 -39
rect 9862 -117 9909 -39
rect 9977 -117 9982 -39
rect 9904 -122 9982 -117
rect 7893 -498 9525 -386
rect 6925 -1593 7052 -1588
rect 6925 -1710 6930 -1593
rect 7047 -1710 7052 -1593
rect 7893 -1610 8005 -498
rect 9413 -728 9525 -498
rect 8289 -840 9525 -728
rect 8289 -1079 8401 -840
rect 8289 -1148 9403 -1079
rect 8289 -1191 9606 -1148
rect 9868 -1186 9933 -1155
rect 6925 -1806 7052 -1710
rect 7888 -1615 8010 -1610
rect 7888 -1717 7893 -1615
rect 8005 -1717 8010 -1615
rect 7888 -1722 8010 -1717
rect 6925 -1931 6926 -1806
rect 7051 -1931 7052 -1806
rect 8344 -1844 8456 -1191
rect 9077 -1260 9606 -1191
rect 9077 -1844 9189 -1260
rect 9494 -1781 9606 -1260
rect 9851 -1677 9963 -1186
rect 10681 -1475 10821 -1470
rect 10681 -1595 10686 -1475
rect 10816 -1595 10821 -1475
rect 10681 -1600 10821 -1595
rect 9851 -1733 9868 -1677
rect 9933 -1733 9963 -1677
rect 9851 -1781 9963 -1733
rect 6926 -1937 7051 -1931
rect 8344 -1956 9224 -1844
rect 9494 -1893 9963 -1781
rect 10686 -1773 10816 -1600
rect 10686 -1907 10816 -1901
rect 9112 -2212 9224 -1956
rect 8404 -2324 9224 -2212
rect 8404 -2516 8516 -2324
rect 7540 -2628 9956 -2516
rect 6927 -3291 7078 -3290
rect 6922 -3296 7083 -3291
rect 6922 -3437 6927 -3296
rect 7078 -3437 7083 -3296
rect 7540 -3437 7652 -2628
rect 7783 -2768 7887 -2652
rect 7944 -2768 8056 -2628
rect 9309 -2661 9389 -2628
rect 7783 -3000 8056 -2768
rect 7783 -3104 7788 -3000
rect 7882 -3104 8056 -3000
rect 7783 -3126 8056 -3104
rect 9290 -2846 9402 -2661
rect 9290 -2916 9309 -2846
rect 9389 -2916 9402 -2846
rect 9290 -3126 9402 -2916
rect 9844 -3126 9956 -2628
rect 7783 -3188 9967 -3126
rect 7783 -3221 7887 -3188
rect 7944 -3238 9967 -3188
rect 6922 -3442 7083 -3437
rect 6927 -3516 7078 -3442
rect 7944 -3456 8056 -3238
rect 9844 -3356 9956 -3238
rect 11097 -3336 11207 -3331
rect 11097 -3426 11102 -3336
rect 11202 -3426 11207 -3336
rect 11097 -3431 11207 -3426
rect 11102 -3506 11202 -3431
rect 11102 -3610 11202 -3604
rect 6927 -3671 7078 -3665
rect 10263 -3729 10408 -3631
rect 11004 -3729 11149 -3725
rect 9923 -3730 11149 -3729
rect 9923 -3762 11009 -3730
rect 8059 -3839 11009 -3762
rect 9923 -3874 11009 -3839
rect 11004 -3875 11009 -3874
rect 11144 -3875 11149 -3730
rect 11004 -3880 11149 -3875
<< via3 >>
rect 8096 -22 8163 43
rect 9786 -117 9862 -39
rect 6926 -1931 7051 -1806
rect 10686 -1901 10816 -1773
rect 6927 -3665 7078 -3516
rect 11102 -3604 11202 -3506
<< metal4 >>
rect 8095 43 8164 44
rect 8095 -22 8096 43
rect 8163 -22 8164 43
rect 8095 -23 8164 -22
rect 8096 -297 8163 -23
rect 9785 -39 9863 -38
rect 9785 -117 9786 -39
rect 9862 -117 9863 -39
rect 9785 -348 9863 -117
rect 9811 -1773 10817 -1772
rect 6925 -1806 7818 -1805
rect 6925 -1931 6926 -1806
rect 7051 -1931 7818 -1806
rect 9811 -1901 10686 -1773
rect 10816 -1901 10817 -1773
rect 9811 -1902 10817 -1901
rect 6925 -1932 7818 -1931
rect 10642 -3506 11203 -3505
rect 6926 -3516 7563 -3515
rect 6926 -3665 6927 -3516
rect 7078 -3665 7563 -3516
rect 10642 -3604 11102 -3506
rect 11202 -3604 11203 -3506
rect 10642 -3605 11203 -3604
rect 6926 -3666 7563 -3665
use JNWTR_CAPX1  JNWTR_CAPX1_0 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 7600 0 1 -1300
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_1
timestamp 1737500400
transform 1 0 9000 0 1 -1300
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_2
timestamp 1737500400
transform 1 0 7600 0 1 -2800
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_3
timestamp 1737500400
transform 1 0 9000 0 1 -2800
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_4
timestamp 1737500400
transform 1 0 7300 0 1 -4200
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_5
timestamp 1737500400
transform 1 0 9700 0 1 -4200
box 0 0 1080 1080
use JNWTR_IVX1_CV  x1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_TR_SKY130A
timestamp 1744212116
transform -1 0 7480 0 -1 -1724
box -150 -120 2130 440
use JNWTR_IVX1_CV  x2
timestamp 1744212116
transform 1 0 10650 0 1 -2080
box -150 -120 2130 440
use JNWTR_IVX1_CV  x12
timestamp 1744212116
transform 1 0 8168 0 1 -4220
box -150 -120 2130 440
use JNWTR_IVX1_CV  x13
timestamp 1744212116
transform -1 0 9886 0 -1 -3300
box -150 -120 2130 440
use JNWATR_NCH_4C5F0  x14 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1744065478
transform 1 0 10384 0 1 -3172
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  x15
timestamp 1744065478
transform 1 0 6234 0 1 -3128
box -184 -128 1336 928
use JNWATR_NCH_2C1F2  xeval1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 8324 0 1 -3032
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch1
timestamp 1734044400
transform -1 0 8508 0 -1 -1051
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch2
timestamp 1734044400
transform 1 0 9144 0 1 -1852
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch3
timestamp 1734044400
transform 1 0 7484 0 1 -1032
box -184 -128 1208 928
use JNWATR_NCH_2C1F2  xlatch4
timestamp 1734044400
transform -1 0 10168 0 -1 -232
box -184 -128 1208 928
use JNWATR_PCH_4C1F2  xpre1 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 5644 0 1 -972
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xpre2
timestamp 1734044400
transform 1 0 5644 0 1 28
box -184 -128 1336 928
use JNWATR_PCH_8C1F2  xpre3 ~/Documents/NTNU/01_Advanced_Integrated_Circuits/aicex/ip/jnw_gr05_sky130a/design/JNW_GR05_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 7104 0 1 28
box -184 -128 1592 928
use JNWATR_PCH_8C1F2  xpre4
timestamp 1734044400
transform -1 0 10552 0 -1 828
box -184 -128 1592 928
use JNWATR_PCH_4C1F2  xpre5
timestamp 1734044400
transform -1 0 12036 0 -1 828
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xpre6
timestamp 1734044400
transform -1 0 12036 0 -1 -172
box -184 -128 1336 928
<< labels >>
flabel metal1 5804 1440 11044 1504 0 FreeSans 1600 0 0 0 CLK
port 6 nsew
flabel metal2 9304 1841 9908 1905 0 FreeSans 1600 0 0 0 Vin2
port 8 nsew
flabel metal2 7790 1841 8284 1905 0 FreeSans 1600 0 0 0 Vin1
port 10 nsew
flabel locali 11358 1012 13366 1204 0 FreeSans 1600 0 0 0 VDD
port 12 nsew
flabel metal1 11056 -3194 12936 -3002 0 FreeSans 1600 0 0 0 Vout
port 14 nsew
flabel locali 10858 -3510 12878 -3318 0 FreeSans 1600 0 0 0 VSS
port 15 nsew
<< properties >>
string FIXED_BBOX 0 0 19740 5720
<< end >>
