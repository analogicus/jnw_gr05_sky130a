* TB_COUNTER_SKY130NM
*----------------------------------------------------------------
* Include Design Files
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_GR05_lpe.spi
#else
.include ../../../work/xsch/JNW_GR05.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param PERIOD_CLK = 100n
.param PW_CLK = {PERIOD_CLK/2}

.param vdda = 1.8
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE (Stimulus)
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  dc {AVDD}

* Clock Source
VCLK clk 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {PW_CLK} {PERIOD_CLK})

* Reset Pulse (Active High)
VRESET reset 0 dc {AVDD} pwl (0 {AVDD} 1n {AVDD} 2n 0)

*-----------------------------------------------------------------
* DUT (Counter)
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi


VB0 b.0 b<0> dc 0
VB1 b.1 b<1> dc 0
VB2 b.2 b<2> dc 0
VB3 b.3 b<3> dc 0
VB4 b.4 b<4> dc 0
*-----------------------------------------------------------------
* PROBES
*-----------------------------------------------------------------
.save all
.save clk reset b[4] b[3] b[2] b[1] b[0]

*----------------------------------------------------------------
* NGSPICE Simulation Control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0

foreach vtemp -20 -10 0 10 20 30 40 50 60 70 80 90 100 110 120
	option temp=$vtemp
	tran 1n 5u 10n
	write {cicname}_$vtemp.raw
end

quit
.endc

.end
